/*
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
NYCU Institute of Electronic
2025 Spring IC Design Laboratory 
Lab09: SystemVerilog Design and Verification 
File Name   : PATTERN.sv
Module Name : PATTERN
Release version : v1.0 (Release Date: April-2025)
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
*/
`define PAT_NUM         8600
`define RANDOM_SEED     5487
// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);
import usertype::*;
//================================================================
// parameters & integer
//================================================================
parameter DRAM_p_r = "../00_TESTBED/DRAM/dram.dat";

parameter MAX_CYCLE=1000;
parameter CLK_TIME = 15;

parameter SEED = `RANDOM_SEED;
integer addr;
integer total_lat, lat;
integer i, i_pat;
//================================================================
// wire & registers 
//================================================================
logic [7:0] golden_DRAM [((65536+8*256)-1):(65536+0)];  // 32 box


Action       action_reg;
Strategy_Type strategy_reg;
Stock stock_A, stock_B, stock_C, stock_D;
Data_No data_reg;
Date date_reg;
Mode         mode_reg;
logic [11:0] Lily_request;
logic [11:0] Rose_request;
logic [11:0] Carnation_request;
logic [11:0] Baby_Breath_request;
logic [63:0] dram_out ,dram_in;
logic overflow_flag;
logic date_check;
logic warn_stock;
Data_Dir dram_in_dir, dram_out_dir;
// Data_Dir dram_in;
Warn_Msg       golden_warn_msg;
logic          golden_complete;
logic [12:0] Lily_new;
logic [12:0] Rose_new;
logic [12:0] Carnation_new;
logic [12:0] Baby_Breath_new;
//================================================================
// class random
//================================================================

/**
 * Class representing a random action.
 */
class random_act;
    randc Action act_id;
    constraint range{
        act_id inside{Purchase, Restock, Check_Valid_Date};
    }
    function new (int seed);
        
        this.srandom(seed);
    endfunction
endclass

class random_strategy;
    randc Strategy_Type strategy_id;
    constraint range{
        strategy_id inside{Strategy_A, Strategy_B, Strategy_C, Strategy_D,
                            Strategy_E, Strategy_F, Strategy_G, Strategy_H};
    }
    function new (int seed);
        
        this.srandom(seed);
    endfunction
endclass

class random_mode;
    randc Mode mode_id;
    constraint range{
        mode_id inside{Single, Group_Order, Event};
    }
    function new(int seed);
        
        this.srandom(seed);
    endfunction
endclass

class random_date;
	randc Date date_id;
	constraint limit{
		date_id.M inside{[1:12]};
        (date_id.M == 1 | date_id.M == 3 | date_id.M == 5 | date_id.M == 7 | date_id.M == 8 | date_id.M == 10 | date_id.M == 12) -> date_id.D inside{[1:31]};
		(date_id.M == 4 | date_id.M == 6 | date_id.M == 9 | date_id.M == 11)                                            -> date_id.D inside{[1:30]};
		(date_id.M == 2)                                                                                       -> date_id.D inside{[1:28]};
	}
    function new(int seed);
        
        this.srandom(seed);
    endfunction
endclass

class random_data_no;
	randc Data_No data_no_id;
	constraint limit{
		data_no_id inside{[0:255]};
	}
    function new(int seed);
        
        this.srandom(seed);
    endfunction
endclass

class random_stock;
    randc Stock stock_id;
    constraint range{
        stock_id inside{[0:4095]};
    }
    function new(int seed);
        
        this.srandom(seed);
    endfunction
endclass
random_act act_rand;
random_strategy strategy_rand;
random_mode mode_rand;
random_date date_rand;
random_data_no data_no_rand;
random_stock stock_rand;
//================================================================
// initial
//================================================================
initial begin
    $readmemh(DRAM_p_r, golden_DRAM);

    act_rand = new(SEED);
    strategy_rand = new(SEED);
    mode_rand = new(SEED);
    date_rand = new(SEED);
    data_no_rand = new(SEED);
    stock_rand = new(SEED);


    reset_task;

    for (i_pat=0; i_pat<`PAT_NUM; i_pat++) begin
        input_task;
        wait_out_valid_task;
        calculate_ans_task;
        $display("inf.warn_msg = %d, inf.complete = %d", inf.warn_msg, inf.complete);
        $display("golden_warn_msg = %d, golden_complete = %d", golden_warn_msg, golden_complete);
        check_ans_task;
		$display("\033[0;34mPASS PATTERN NO.%4d, \033[m \033[0;32m Execution Cycle: %3d\033[m", i_pat, lat);
    end
    YOU_PASS_task;
    $finish;
end



//================================================================
// task
//================================================================
task reset_task; begin
    inf.rst_n = 1'b1;

    inf.sel_action_valid = 1'b0;
    inf.strategy_valid = 1'b0;
    inf.mode_valid = 1'b0;
    inf.date_valid = 1'b0;
    inf.data_no_valid = 1'b0;
    inf.restock_valid = 1'b0;
    inf.D = 'dx;

    #(1); inf.rst_n = 0;
    #(5); inf.rst_n = 1;
end
endtask


task input_task; begin
    @(negedge clk);
    inf.sel_action_valid = 1;
    act_rand.randomize();
    action_reg = act_rand.act_id;
    inf.D.d_act[0] = action_reg; 
    @(negedge clk); 
	inf.sel_action_valid = 0; 
    inf.D = 'bx;

    case (action_reg)
        Purchase: begin
            repeat($urandom_range(0,3))@(negedge clk);
            input_strategy_task;
            repeat($urandom_range(0,3))@(negedge clk);
            input_mode_task;
            repeat($urandom_range(0,3))@(negedge clk);
            input_date_task;
            repeat($urandom_range(0,3))@(negedge clk);
            input_data_no_task;
        end
        Restock: begin
            repeat($urandom_range(0,3))@(negedge clk);
            input_date_task;
            repeat($urandom_range(0,3))@(negedge clk);
            input_data_no_task;
            input_restock_task;
        end
        Check_Valid_Date: begin
            repeat($urandom_range(0,3))@(negedge clk);
            input_date_task;
            repeat($urandom_range(0,3))@(negedge clk);
            input_data_no_task;
        end
    endcase
end
endtask

task input_strategy_task; begin
    inf.strategy_valid = 1'd1;
    strategy_rand.randomize();
    strategy_reg = strategy_rand.strategy_id;
    inf.D.d_strategy[0] = strategy_reg;
    @(negedge clk); 
    inf.strategy_valid = 1'd0;
    inf.D = 'bx;
end
endtask
task input_mode_task; begin
    inf.mode_valid = 1'd1;
    mode_rand.randomize();
    mode_reg = mode_rand.mode_id;
    inf.D.d_mode[0] = mode_reg;
    @(negedge clk); 
    inf.mode_valid = 1'd0;
    inf.D = 'bx;
end
endtask
task input_date_task; begin
    inf.date_valid = 1'd1;
    date_rand.randomize();
    date_reg = date_rand.date_id;
    inf.D.d_date[0] = date_reg;
    @(negedge clk); 
    inf.date_valid = 1'd0;
    inf.D = 'bx;
end
endtask
task input_data_no_task; begin
    inf.data_no_valid = 1'd1;
    data_no_rand.randomize();
    data_reg = data_no_rand.data_no_id;
    inf.D.d_data_no[0] = data_reg;
    @(negedge clk); 
    inf.data_no_valid = 1'd0;
    inf.D = 'bx;
end
endtask

task input_restock_task; begin
    for (i = 0 ; i < 4 ; i++) begin
        repeat($urandom_range(0,3))@(negedge clk);
        inf.restock_valid = 1'd1;
        stock_rand.randomize();
        inf.D.d_stock[0]= stock_rand.stock_id;
        case (i)
            0    : stock_A = inf.D.d_stock[0];
            1    : stock_B = inf.D.d_stock[0];
            2    : stock_C = inf.D.d_stock[0];
            3    : stock_D = inf.D.d_stock[0]; 
        endcase
        @(negedge clk); 
        inf.restock_valid = 1'd0;
        inf.D = 'bx;
    end
end
endtask

task wait_out_valid_task; begin
  lat = -1; 
  while(inf.out_valid !== 1) begin 
  	lat = lat + 1;  
		if(lat == 1000) begin
            YOU_FAIL_task;
            $display("--------------------------------------------------------------------------------------------------------------------------------------------");
            $display("                                                             PATTERN NO.%4d 	                                                              ", i_pat);
            $display("                                             The execution latency should not over 1000 cycles                                              ");
            $display("--------------------------------------------------------------------------------------------------------------------------------------------");
            $finish;
		end
	@(negedge clk);
  end
  total_lat = total_lat + lat;
end
endtask


task calculate_ans_task; begin
    addr = 65536 + 8 * data_reg;
     dram_out = {golden_DRAM[addr+7], golden_DRAM[addr+6], golden_DRAM[addr+5], golden_DRAM[addr+4], golden_DRAM[addr+3], golden_DRAM[addr+2], golden_DRAM[addr+1], golden_DRAM[addr]};
     dram_out_dir.Rose       = dram_out[63:52];
     dram_out_dir.Lily       = dram_out[51:40];
     dram_out_dir.M          = dram_out[39:32];
     dram_out_dir.Carnation  = dram_out[31:20];
     dram_out_dir.Baby_Breath= dram_out[19:8];
     dram_out_dir.D          = dram_out[7:0];

    $display("DEBUG: action_reg = %0d", action_reg);
    $display("DEBUG: data_reg = %0d", data_reg);
    $display("DEBUG: date_reg.M = %0d", date_reg.M);
    $display("DEBUG: date_reg.D = %0d", date_reg.D);
    $display("DEBUG: strategy_reg = %0d, mode_reg = %0d", strategy_reg, mode_reg);
    $display("DEBUG: After all cases, dram_out_dir.Rose = %0d", dram_out_dir.Rose);
    $display("DEBUG: After all cases, dram_out_dir.Lily = %0d", dram_out_dir.Lily);
    $display("DEBUG: After all cases, dram_out_dir.M = %0d", dram_out_dir.M);
    $display("DEBUG: After all cases, dram_out_dir.D = %0d", dram_out_dir.D);
    $display("DEBUG: After all cases, dram_out_dir.Carnation = %0d", dram_out_dir.Carnation);
    $display("DEBUG: After all cases, dram_out_dir.Baby_Breath = %0d", dram_out_dir.Baby_Breath);
    // date_check = (date_reg.M < dram_out_dir.M) | ((date_reg.M == dram_out_dir.M) & (date_reg.D < dram_out_dir.D)) && action_reg != Restock  ;
    // overflow_flag = Lily_new[12] | Rose_new[12] | Carnation_new[12] | Baby_Breath_new[12];
    // warn_stock = ( (dram_out_dir.Rose < Rose_request) | (dram_out_dir.Lily < Lily_request) | (dram_out_dir.Carnation < Carnation_request) | (dram_out_dir.Baby_Breath < Baby_Breath_request));

    if (action_reg == Purchase) begin
        // $display("DEBUG: In Purchase case, strategy_reg = %0d, mode_reg = %0d", strategy_reg, mode_reg);
        Lily_request = 0;
        Rose_request = 0;
        Carnation_request = 0;
        Baby_Breath_request = 0;
         case (strategy_reg)
            Strategy_A: begin
                case (mode_reg)
                    Single: begin
                        Rose_request = 'd120;
                        // $display("DEBUG: In Single mode case, setting Rose_request to 120");
                    end
                    Group_Order: begin
                        Rose_request = 'd480;
                    end
                    Event: begin
                        Rose_request = 'd960;
                    end
                    default: begin
                        Rose_request = 0;
                    end
                endcase
            end
            Strategy_B: begin
                case (mode_reg)
                    Single: begin
                        Lily_request = 'd120;
                    end
                    Group_Order: begin
                        Lily_request = 'd480;
                    end
                    Event: begin
                        Lily_request = 'd960;
                    end
                    default: begin
                        Lily_request = 0;
                    end
                endcase
            end
            Strategy_C: begin
                case (mode_reg)
                    Single: begin
                        Carnation_request = 'd120;
                    end
                    Group_Order: begin
                        Carnation_request = 'd480;
                    end
                    Event: begin
                        Carnation_request = 'd960;
                    end
                    default: begin
                        Carnation_request = 0;
                    end
                endcase
            end
            Strategy_D: begin
                case (mode_reg)
                    Single: begin
                        Baby_Breath_request = 'd120;
                    end
                    Group_Order: begin
                        Baby_Breath_request = 'd480;
                    end
                    Event: begin
                        Baby_Breath_request = 'd960;
                    end
                    default: begin
                        Baby_Breath_request = 0;
                    end
                endcase
            end
            Strategy_E: begin
                case (mode_reg)
                    Single: begin
                        Rose_request = 'd60;
                        Lily_request = 'd60;
                    end
                    Group_Order: begin
                        Rose_request = 'd240;
                        Lily_request = 'd240;
                    end
                    Event: begin
                        Rose_request = 'd480;
                        Lily_request = 'd480;
                    end
                    default: begin
                        Rose_request = 'd0;
                        Lily_request = 'd0;
                    end
                endcase
            end
            Strategy_F: begin
                case (mode_reg)
                    Single: begin
                        Carnation_request = 'd60;
                        Baby_Breath_request = 'd60;
                    end
                    Group_Order: begin
                        Carnation_request = 'd240;
                        Baby_Breath_request = 'd240;
                    end
                    Event: begin
                        Carnation_request = 'd480;
                        Baby_Breath_request = 'd480;
                    end
                    default: begin
                        Carnation_request = 'd0;
                        Baby_Breath_request = 'd0;
                    end
                endcase
            end
            Strategy_G: begin
                case (mode_reg)
                    Single: begin
                        Carnation_request = 'd60;
                        Rose_request = 'd60;
                    end
                    Group_Order: begin
                        Carnation_request = 'd240;
                        Rose_request = 'd240;
                    end
                    Event: begin
                        Carnation_request = 'd480;
                        Rose_request = 'd480;
                    end
                    default: begin
                        Carnation_request = 'd0;
                        Rose_request = 'd0;
                    end
                endcase
            end
            Strategy_H: begin
                case (mode_reg)
                    Single: begin
                        Carnation_request = 'd30;
                        Baby_Breath_request = 'd30;
                        Rose_request = 'd30;
                        Lily_request = 'd30;
                    end
                    Group_Order: begin
                        Carnation_request = 'd120;
                        Baby_Breath_request = 'd120;
                        Rose_request = 'd120;
                        Lily_request = 'd120;
                    end
                    Event: begin
                        Carnation_request = 'd240;
                        Baby_Breath_request = 'd240;
                        Rose_request = 'd240;
                        Lily_request = 'd240;
                    end
                    default: begin
                        Carnation_request = 'd0;
                        Baby_Breath_request = 'd0;
                        Rose_request = 'd0;
                        Lily_request = 'd0;
                    end
                endcase
            end 
         endcase
         $display("DEBUG: After all cases, Rose_request = %0d", Rose_request);
         $display("DEBUG: After all cases, Lily_request = %0d", Lily_request);
         $display("DEBUG: After all cases, Carnation_request = %0d", Carnation_request);
         $display("DEBUG: After all cases, Baby_Breath_request = %0d", Baby_Breath_request);
        //  $display("DEBUG: After all cases, dram_out_dir.Rose = %0d", dram_out_dir.Rose);
        //  $display("DEBUG: After all cases, dram_out_dir.Lily = %0d", dram_out_dir.Lily);
        //  $display("DEBUG: After all cases, dram_out_dir.Carnation = %0d", dram_out_dir.Carnation);
        //  $display("DEBUG: After all cases, dram_out_dir.Baby_Breath = %0d", dram_out_dir.Baby_Breath);
        //  if (( (dram_out_dir.Rose < Rose_request) || (dram_out_dir.Lily < Lily_request) || (dram_out_dir.Carnation < Carnation_request) || (dram_out_dir.Baby_Breath < Baby_Breath_request))) begin
        //     golden_complete = 0;
        //     golden_warn_msg = Stock_Warn;
        //  end
         if ((date_reg.M < dram_out_dir.M) || ((date_reg.M == dram_out_dir.M) && (date_reg.D < dram_out_dir.D)))  begin
            golden_complete = 0;
            golden_warn_msg = Date_Warn;
         end
         else if (( (dram_out_dir.Rose < Rose_request) || (dram_out_dir.Lily < Lily_request) || (dram_out_dir.Carnation < Carnation_request) || (dram_out_dir.Baby_Breath < Baby_Breath_request))) begin
            golden_complete = 0;
            golden_warn_msg = Stock_Warn;
         end
        //  if (!(date_reg.M < dram_out_dir.M) || ((date_reg.M == dram_out_dir.M) && (date_reg.D < dram_out_dir.D)) && !( (dram_out_dir.Rose < Rose_request) | (dram_out_dir.Lily < Lily_request) | (dram_out_dir.Carnation < Carnation_request) | (dram_out_dir.Baby_Breath < Baby_Breath_request))) 
         else
         begin
            golden_complete = 1;
            golden_warn_msg = No_Warn;
            dram_in_dir.Rose       = dram_out_dir.Rose - Rose_request;
            dram_in_dir.Lily       = dram_out_dir.Lily - Lily_request;
            dram_in_dir.Carnation  = dram_out_dir.Carnation - Carnation_request;
            dram_in_dir.Baby_Breath= dram_out_dir.Baby_Breath - Baby_Breath_request;
            dram_in_dir.M          = dram_out_dir.M;
            dram_in_dir.D          = dram_out_dir.D;
            dram_in = {dram_in_dir.Rose, dram_in_dir.Lily,4'b0000 ,dram_in_dir.M, dram_in_dir.Carnation, dram_in_dir.Baby_Breath,3'b000 ,dram_in_dir.D};
            {golden_DRAM[addr+7], golden_DRAM[addr+6], golden_DRAM[addr+5], golden_DRAM[addr+4], golden_DRAM[addr+3], golden_DRAM[addr+2], golden_DRAM[addr+1], golden_DRAM[addr]} = dram_in;
         end
    end else if (action_reg == Restock) begin
        // calculate ans for Restock action
        golden_complete = 1;
        golden_warn_msg = No_Warn;
        
        Lily_new = dram_out_dir.Lily + stock_B;
        Rose_new = dram_out_dir.Rose + stock_A;
        Carnation_new = dram_out_dir.Carnation + stock_C;
        Baby_Breath_new = dram_out_dir.Baby_Breath + stock_D;
        if (Lily_new[12] || Rose_new[12] || Carnation_new[12] || Baby_Breath_new[12]) begin
            golden_complete = 0;
            golden_warn_msg = Restock_Warn;
        end
        dram_in_dir.M           = date_reg.M;
        dram_in_dir.D           = date_reg.D;
        dram_in_dir.Lily        = Lily_new[12]==1        ? 12'd4095 : Lily_new[11:0];
        dram_in_dir.Rose        = Rose_new[12]==1        ? 12'd4095 : Rose_new[11:0];
        dram_in_dir.Carnation   = Carnation_new[12]==1   ? 12'd4095 : Carnation_new[11:0];
        dram_in_dir.Baby_Breath = Baby_Breath_new[12]==1 ? 12'd4095 : Baby_Breath_new[11:0];
        dram_in = {dram_in_dir.Rose, dram_in_dir.Lily,4'b0000 ,dram_in_dir.M, dram_in_dir.Carnation, dram_in_dir.Baby_Breath,3'b000 ,dram_in_dir.D};
        {golden_DRAM[addr+7], golden_DRAM[addr+6], golden_DRAM[addr+5], golden_DRAM[addr+4], golden_DRAM[addr+3], golden_DRAM[addr+2], golden_DRAM[addr+1], golden_DRAM[addr]} = dram_in;
    end else if (action_reg == Check_Valid_Date) begin
        // calculate ans for Check_Valid_Date action
        if ((date_reg.M < dram_out_dir.M) || ((date_reg.M == dram_out_dir.M) && (date_reg.D < dram_out_dir.D))) begin
            golden_complete = 0;
            golden_warn_msg = Date_Warn;
        end else begin
            golden_complete = 1;
            golden_warn_msg = No_Warn;
        end
    end 
end
    $display("DEBUG: After all cases, dram_in_dir.Rose = %0d", dram_in_dir.Rose);
    $display("DEBUG: After all cases, dram_in_dir.Lily = %0d", dram_in_dir.Lily);
    $display("DEBUG: After all cases, dram_in_dir.M = %0d", dram_in_dir.M);
    $display("DEBUG: After all cases, dram_in_dir.D = %0d", dram_in_dir.D);
    $display("DEBUG: After all cases, dram_in_dir.Carnation = %0d", dram_in_dir.Carnation);
    $display("DEBUG: After all cases, dram_in_dir.Baby_Breath = %0d", dram_in_dir.Baby_Breath);
endtask

// task check_ans_task; begin
//     if((inf.warn_msg !== golden_warn_msg) | (inf.complete !== golden_complete)) begin
//         $display(" \033[0;31m ");
//         $display(" Wrong Answer ");
//         $display(" \033[m ");
//         $finish;
//     end
// end endtask

task check_ans_task; begin
   if(inf.out_valid ===1) begin 
    if((inf.complete !== golden_complete) || (inf.warn_msg !== golden_warn_msg)) begin
        $display("--------------------------------------------------------------------------------------------------------------------------------------------");
        $display("                                                             PATTERN NO.%4d 	                                                              ", i_pat);
        $display("                                             The output complete is wrong, please check it!                                              ");
        $display("--------------------------------------------------------------------------------------------------------------------------------------------");
        $finish;
    end
    // if(inf.warn_msg !== golden_warn_msg) begin
    //     $display("--------------------------------------------------------------------------------------------------------------------------------------------");
    //     $display("                                                             PATTERN NO.%4d 	                                                              ", i_pat);
    //     $display("                                             The output warn_msg is wrong, please check it!                                              ");
    //     $display("--------------------------------------------------------------------------------------------------------------------------------------------");
    //     $finish;
    // end
    
   end
@(negedge inf.out_valid);

end endtask




task YOU_PASS_task; begin
	$display("\033[37m                                  .$&X.      x$$x              \033[32m      :BBQvi.");
	$display("\033[37m                                .&&;.X&$  :&&$+X&&x            \033[32m     BBBBBBBBQi");
	$display("\033[37m                               +&&    &&.:&$    .&&            \033[32m    :BBBP :7BBBB.");
	$display("\033[37m                              :&&     &&X&&      $&;           \033[32m    BBBB     BBBB");
	$display("\033[37m                              &&;..   &&&&+.     +&+           \033[32m   iBBBv     BBBB       vBr");
	$display("\033[37m                             ;&&...   X&&&...    +&.           \033[32m   BBBBBKrirBBBB.     :BBBBBB:");
	$display("\033[37m                             x&$..    $&&X...    +&            \033[32m  rBBBBBBBBBBBR.    .BBBM:BBB");
	$display("\033[37m                             X&;...   &&&....    &&            \033[32m  BBBB   .::.      EBBBi :BBU");
	$display("\033[37m                             $&...    &&&....    &&            \033[32m MBBBr           vBBBu   BBB.");
	$display("\033[37m                             $&....   &&&...     &$            \033[32m i7PB          iBBBBB.  iBBB");
	$display("\033[37m                             $&....   &&& ..    .&x                        \033[32m  vBBBBPBBBBPBBB7       .7QBB5i");
	$display("\033[37m                             $&....   &&& ..    x&+                        \033[32m :RBBB.  .rBBBBB.      rBBBBBBBB7");
	$display("\033[37m                             X&;...   x&&....   &&;                        \033[32m    .       BBBB       BBBB  :BBBB");
	$display("\033[37m                             x&X...    &&....   &&:                        \033[32m           rBBBr       BBBB    BBBU");
	$display("\033[37m                             :&$...    &&+...   &&:                        \033[32m           vBBB        .BBBB   :7i.");
	$display("\033[37m                              &&;...   &&$...   &&:                        \033[32m             .7  BBB7   iBBBg");
	$display("\033[37m                               && ...  X&&...   &&;                                         \033[32mdBBB.   5BBBr");
	$display("\033[37m                               .&&;..  ;&&x.    $&;.$&$x;                                   \033[32m ZBBBr  EBBBv     YBBBBQi");
	$display("\033[37m                               ;&&&+   .+xx;    ..  :+x&&&&&&&x                             \033[32m  iBBBBBBBBD     BBBBBBBBB.");
	$display("\033[37m                        +&&&&&&X;..             .          .X&&&&&x                         \033[32m    :LBBBr      vBBBi  5BBB");
	$display("\033[37m                    $&&&+..                                    .:$&&&&.                     \033[32m          ...   :BBB:   BBBu");
	$display("\033[37m                 $&&$.                                             .X&&&&.                  \033[32m         .BBBi   BBBB   iMBu");
	$display("\033[37m              ;&&&:                                               .   .$&&&                x\033[32m          BBBX   :BBBr");
	$display("\033[37m            x&&x.      .+&&&&&.                .x&$x+:                  .$&&X         $+  &x  ;&X   \033[32m  .BBBv  :BBBQ");
	$display("\033[37m          .&&;       .&&&:                      .:x$&&&&X                 .&&&        ;&     +&.    \033[32m   .BBBBBBBBB:");
	$display("\033[37m         $&&       .&&$.                             ..&&&$                 x&& x&&&X+.          X&x\033[32m     rBBBBB1.");
	$display("\033[37m        &&X       ;&&:                                   $&&x                $&x   .;x&&&&:                       ");
	$display("\033[37m      .&&;       ;&x                                      .&&&                &&:       .$&&$    ;&&.             ");
	$display("\033[37m      &&;       .&X                                         &&&.              :&$          $&&x                   ");
	$display("\033[37m     x&X       .X& .                                         &&&.              .            ;&&&  &&:             ");
	$display("\033[37m     &&         $x                                            &&.                            .&&&                 ");
	$display("\033[37m    :&&                                                       ;:                              :&&X                ");
	$display("\033[37m    x&X                 :&&&&&;                ;$&&X:                                          :&&.               ");
	$display("\033[37m    X&x .              :&&&  $&X              &&&  X&$                                          X&&               ");
	$display("\033[37m    x&X                x&&&&&&&$             :&&&&$&&&                                          .&&.              ");
	$display("\033[37m    .&&    \033[38;2;255;192;203m      ....\033[37m  .&&X:;&&+              &&&++;&&                                          .&&               ");
	$display("\033[37m     &&    \033[38;2;255;192;203m  .$&.x+..:\033[37m  ..+Xx.                 :&&&&+\033[38;2;255;192;203m  .;......    \033[37m                             .&&");
	$display("\033[37m     x&x   \033[38;2;255;192;203m .x&:;&x:&X&&.\033[37m              .             \033[38;2;255;192;203m .&X:&&.&&.:&.\033[37m                             :&&");
	$display("\033[37m     .&&:  \033[38;2;255;192;203m  x;.+X..+.;:.\033[37m         ..  &&.            \033[38;2;255;192;203m &X.;&:+&$ &&.\033[37m                             x&;");
	$display("\033[37m      :&&. \033[38;2;255;192;203m    .......   \033[37m         x&&&&&$++&$        \033[38;2;255;192;203m .... ......: \033[37m                             && ");
	$display("\033[37m       ;&&                          X&  .x.              \033[38;2;255;192;203m .... \033[37m                               .&&;                ");
	$display("\033[37m        .&&x                        .&&$X                                          ..         .x&&&               ");
	$display("\033[37m          x&&x..                                                                 :&&&&&+         +&X              ");
	$display("\033[37m            ;&&&:                                                                     x&&$XX;::x&&X               ");
	$display("\033[37m               &&&&&:.                                                              .X&x    +xx:                  ");
	$display("\033[37m                  ;&&&&&&&&$+.                                  :+x&$$X$&&&&&&&&&&&&&$                            ");
	$display("\033[37m                       .+X$&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&$X+xXXXxxxx+;.                                   ");
end endtask

task YOU_FAIL_task; begin                                                                                                                         
	$display("\033[37m                                                                         x&&&&X  +&&&&&&+                                    ");
	$display("\033[37m                                                                      .&&&&$$&&&&&&+ .&&&&                                   ");
	$display("\033[37m                                                                     X&&&;   &&&&$     X&&&                                  ");
	$display("\033[31m i:..::::::i.      :::::         ::::    .:::.        \033[37m              &&&X.    &&&&..    .&&&;                                 ");
	$display("\033[31m BBBBBBBBBBBi     iBBBBBL       .BBBB    7BBB7        \033[37m             &&&X .   .&&&; .    .&&&;                                 ");
	$display("\033[31m BBBB.::::ir.     BBB:BBB.      .BBBv    iBBB:        \033[37m            X&&&...   +&&&. .    ;&&&:                                 ");
	$display("\033[31m BBBQ            :BBY iBB7       BBB7    :BBB:        \033[37m           ;&&&; ..  .&&&X  .    x&&&.                                 ");
	$display("\033[31m BBBB            BBB. .BBB.      BBB7    :BBB:        \033[37m           &&&$  ..  ;&&&+  .   .&&&$                                  ");
	$display("\033[31m BBBB:r7vvj:    :BBB   gBBs      BBB7    :BBB:        \033[37m          .&&&;  ..  $&&&. ..   ;&&&;                                  ");
	$display("\033[31m BBBBBBBBBB7    BBB:   .BBB.     BBB7    :BBB:        \033[37m          ;&&&:  .  .&&&x ..    X&&&                                   ");
	$display("\033[31m BBBB    ..    iBBBBBBBBBBBP     BBB7    :BBB:        \033[37m          +&&&.  .  +&&&: ..   .&&&x                                   ");
	$display("\033[31m BBBB          BBBBi7vviQBBB.    BBB7    :BBB.        \033[37m          +&&&.     $&&X. ..   X&&&.                                   ");
	$display("\033[31m BBBB         rBBB.      BBBQ   .BBBv    iBBB2ir777L7 \033[37m          +&&&.    :&&&:...   :&&&X                                    ");
	$display("\033[31m.BBBB        :BBBB       BBBB7  .BBBB    7BBBBBBBBBBB \033[37m          ;&&&.    x&&$       X&&&.                                    ");
	$display("\033[31m . ..        ....         ...:   ....    ..   ....... \033[37m          .&&&.   .&&&&+.    :&&&X                                     ");
	$display("\033[37m                                                        :+X&&.   X&X     X&&&X.    &&&&                                      ");
	$display("\033[37m                                                    ;$&&&&&&&:                     :Xx  ;&&&&&&$;                            ");
	$display("\033[37m                                                .$&&&&&X;.                                 ;x&&&&&&+   $&&&X:                ");
	$display("\033[37m                                              ;&&&&&x.                                         :$&&&&;  ;x&&&&&:             ");
	$display("\033[37m                                            :&&&&&.      .;X$$:                   ....            ;&&&&+    .x&&&x           ");
	$display("\033[37m                                           $&&&x.     .$&&&&&&x.                ;&&&&&&&$;          :&&&&;      $&&X         ");
	$display("\033[37m                                         :&&&&.     .$&&&;.                        ..;&&&&&$.         x&&&x      :&&&.       ");
	$display("\033[37m                                        .&&&&      :&&&.                                ;&&&&:         +&&&x       $&&+      ");
	$display("\033[37m                                        $&&$.     :&&X                                   .$&&&:         ;&&&+       &&&x     ");
	$display("\033[37m                                       x&&&.     .&&x                                   .  &&&&.         $&&&:      .&&&+    ");
	$display("\033[37m                                      :&&&:       ;+.      .:;:..              :&&&&&x     :&&&.         ;&&&x       +&&&    ");
	$display("\033[37m                                      X&&$               .&&&&&&&&.           X&&& .&&&+     .           .&&&$       :&&&;   ");
	$display("\033[37m                                      &&&;               $&&& +&&&X           $&&&&&&&&x                  $&&&:       &&&&   ");
	$display("\033[37m                                     +&&&.               X&&&&&&&&;           +&&&&x&&&.             .    x&&&;       x&&&:  ");
	$display("\033[37m                                     &&&X  \033[38;2;255;192;203m      ....   \033[37m .X&&&&&&;             .x&&&&X.\033[38;2;255;192;203m  ......    \033[37m  ..   ;&&&:       +&&&+  ");
	$display("\033[37m                                     X&&X  \033[38;2;255;192;203m  .  ;&$. .. \033[37m                .              \033[38;2;255;192;203m x&&:   ..  \033[37m       +&&&.       ;&&&+  ");
	$display("\033[37m         x&&&&&&&&&&&&&&&&&X         +&&$  \033[38;2;255;192;203m .. .&&&:&&&: . \033[37m        .:..&&&;          \033[38;2;255;192;203m .+&&&.x&&: . \033[37m       x&&&        :&&&X  ");
	$display("\033[37m      :;  xxxx;   .;;;.  .$&&.       :&&&. \033[38;2;255;192;203m  . .XX.x&&;  . \033[37m       .&&&&&&&&&X;       \033[38;2;255;192;203m ..&&:.$&&&.. \033[37m      .&&&X        ;&&&x  ");
	$display("\033[37m   ;&&&&:                  x&&:       $&&$ \033[38;2;255;192;203m        .:.. .  \033[37m         +&&&;x&&&x.      \033[38;2;255;192;203m .      .:.   \033[37m      ;&&&.        ;&&&;  ");
	$display("\033[37m :&&&&&&$        .+$&&&$Xx+X&&&.       &&&X\033[38;2;255;192;203m    ........    \033[37m         .&&&+            \033[38;2;255;192;203m    .......   \033[37m     .&&&x         X&&&   ");
	$display("\033[37m &&$   +&&&&&&&&&&&&&&&&&&&&&&&;       .&&&&.                        ;&&&&.                             X&&&          &&&$   ");
	$display("\033[37m &&x:&x  $&&&&&&X.          x&&         .&&&&+                         .:.                             X&&&          .&&&;   ");
	$display("\033[37m.&&$:&&+ :&&;x&&            $&&           :&&&&;                                                     ;&&&X           x&&&    ");
	$display("\033[37m X&&&:   .&&; &&+           ;&&;             $&&$.                                                  ;&&&             &&&+    ");
	$display("\033[37m  :&&&&$$&&&&$&&&            $&&.            ;&&+                                                    .&&;           x&&&.    ");
	$display("\033[37m     x&&&&&&&&&&&;           x&&&+           $&&.     .                                   ;&&+       .&&X          :&&&+     ");
	$display("\033[37m               +&&. .+x$&&&&&&&X:            &&&.   .&&$                                 x&&X  .&$   .&&X         +&&&;      ");
	$display("\033[37m                &&&&&&&&&&&X:                &&&.   .&&;                                .&&&+ ;&&&.  ;&&&+        &&$        ");
	$display("\033[37m                 ;+:                         +&&$. +&&X                                  $&&&&&&&;   X&&&&X                  ");
	$display("\033[37m                                              :&&&&&&&+.                                 .+&&&&;    :&&&&&&.   :&$           ");
	$display("\033[37m                                                     &&&;                                          .&&&&&&&    X&&+          ");
	$display("\033[37m                                                     .&&&:                                        .&&&&&&&     &&&&          ");
	$display("\033[37m                                                      :&&&;                                      ;&&&&&&&x    x&&&x          ");
	$display("\033[37m                                                   :&x  &&&$.                                   x&&&&&&&.    $&&&&$          ");
	$display("\033[37m                                                  +&&X    x&&&&;                              x&&&&&&&x    .&&&&&&&          ");
	$display("\033[37m                                                  &&&       x&&+    +$;      ..        ..;X&&&&&&&&x.     x&&&&&&&X          ");
	$display("\033[37m                                                  $&&       .&&&   :&&&.   .$&&:&&&&&&&&&&&&&$;          &&&&X &&&;          ");
	$display("\033[37m                                                  :&&&:      +&&&;;&&&&    X&&. x&&&&&$X:             .$&&&&: ;&&&           ");
	$display("\033[37m                                                   ;&&&$      .$&&&&&&&$:X&&$                       :&&&&&:  :&&&:           ");
	$display("\033[37m                                                    .&&&&&;          X&&&&X.                     +&&&&&X    +&&&.            ");
	$display("\033[37m                                                      .$&&&&&+                               x&&&&&&+      ;&&&.             ");
	$display("\033[37m                                                         :&&&&&&&&$+.            .;+xX$&&&&&&&&&X:        +&&&:              ");
	$display("\033[37m                                                           $&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&x:           +&&&&.               ");
	$display("\033[37m                                                             x&&&&;+X&&&&&&&&&&&$x.                  :$&&&&:                 ");
	$display("\033[37m                                                               &&&&$:                             .X&&&&x                    ");
	$display("\033[37m                                                                .&&&&&&&&&&+                   X&&&&&$.                      ");
	$display("\033[37m                                                                      .;&&&&&                  $&&&+                         ");
	$display("\033[37m                                                                         &&&&+.             :x&&&&:                          ");
	$display("\033[37m                                                                          X&&&&&&&&&&&&&&&&&&&&$                             ");
	$display("\033[37m                                                                             .;xX$&&&&&$$x+:                                 ");
end endtask
endprogram








/*
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
NYCU Institute of Electronic
2025 Spring IC Design Laboratory 
Lab09: SystemVerilog Design and Verification 
File Name   : PATTERN.sv
Module Name : PATTERN
Release version : v1.0 (Release Date: April-2025)
//   (C) Copyright Laboratory System Integration and Silicon Implementation
//   All Right Reserved
++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++
*/
// `include "../00_TESTBED/pseudo_DRAM.sv"

// `define PAT_NUM     10000
// `define SEED        5487

// `include "Usertype.sv"

// program automatic PATTERN(input clk, INF.PATTERN inf);

// `protected
// 7IO<O>Fd8gFE_&Y>JDe?dHUc9[=b2aO4,FLR>DFd->53G+6=3>X#3)[]4a7[Z8WG
// 6CfbgVUZKAaAYXUA#=LC?+ff83a7)PP5V?N.BNOEc+HHd>.@5H6aYDBQW74.H19A
// 9<4C_<.Y:Q9O]99T+[8e>)+#ZL3NM#aggccM]I=L3JcV>BM80(3:L[CgcS6Kf[Vg
// /WIHMe^OW9]6/TXfB2HH@?C;M+<(,?SIC,/+;TPad;+&G7L&M#(<G;6M(M]^e\.^
// 4aWS?bA2KHT^N]Y)eQ:DcYH,2.Y:/F0BE.3B:P\@8]5S;O03+0aK3NQgNX&D^_]J
// LJ/Ddcgf>d3\^]FI@8C9IaYMc_W#&gO/=OBWP0@aA.?Y]8JN3RM&Vb#D>TCB3bK4
// \d19,]FN[8_aB&T8B/?HZQX=[O2CN.8?8d6eK_W85J5B;eS4(GULd=A+Y926;KE7
// G(RbW3I+#gN&2X#WRHWJcGYVWT+U,e7NJ@:,aD6;-@V6.eTHAA@<0-O+S/3KDY^O
// fTD_<S44g]X4ReT7NB(3GWgVPQ4>bXaWGT3RK;2dD9W?(;1WN4R/;PVBC<#+cWJU
// W5EXX-aMQE^84@3MJ61]]#)\\9V<>R)_e4+@McTJ@_278^a/c]H[bA-]5974Led;
// 4Jdb-aWDOEQ::Z]Q<]_T\A<eN_D5J^XY([ZG;>;-E)1\K49Z,[,T3+8<cTBf\b]5
// +00Ge\5=AUZHdb<]_T;3^3dRN4Q=VZFUdYP6+.[IV-caW+JW?Xa23YOM_VZHW?N=
// [RP&^&U^d2;Ge2GADC]4)_f:g=OX/)HM;SD0NEK1Y.^C<+bG,6O-TD<fRSXTGE6U
// \G6&f?X\,JYgH)FIN7f_S?9Sg10ROBUb&IMU#Q/?#ZK20,\(L)ZLWDb3XJ2,<7B]
// 9fOBXQBZ]fP0:P<R;&2S5Y(Z@F4RI@-P?<NMa52^.QdIdXRO#Q+D^\Vc-Sb)a>;.
// >]TbP3f=-a,eP05Z6RQMHY<#N@TIPf7^9:&GbY]VU/D1Yf_2C\Ve9+Ve#UC5D&Y.
// .E9B_OBdE]0C&2]Q93Me8=dU7;<+HDWKIY(eMZ[6XM59PA)&([O@SG>HP5f(cLD]
// Vef##6\T?].P1Sg[IJLP5&8\?c[,:BMV[CA25NH[eDG/RUS1.fM7M0S+,K167b-F
// E6IA95B+ACTXd4AM-#,KIe2;T>d1THeU?bTb>@fYdDKF2IJLdX6f@d8S4[)6;<;Z
// WEb^-^Yf\C]BYZHH^-)F44\WCP&H5dR=7M5eB@/].=YX+>XJV<Z.4IF\Z.^N_@:I
// ,a<<0?4X(=/.G[I:D?2&4dXPC+CJ@aLLG(MbSZ#cX83^I0BXX?77J<?AA=_MM+5E
// g0=Q)P[92KQ:QG&JUCfVME);FD&4=5)#7cPPg9N-E7GFG]g1H];a(>99[7c71P>9
// 3&d+9,H074U/[O)FTD8GK2],G,1R<S6)^YW6_]S8>:C5ND1Abc37@8M@gd5?0:NN
// 3ZG:09BB[WR\^Rc=(gD/D15XA&-&TdX@KV=I@NVc:_I\7Q5JXbA>F?UbKG,>O[/?
// NID2\EK(/AS6ZWd8PDZ>X6>1SEI#56P^ZJWdc=f4.^85b0(.BTR&N>K5CFH7JETI
// &R3CbE[<H6]>3BV\W,>b;.?+-gXE9?@K/cbcUS.RPJ37C18;A/GdN:](+Je5cZKg
// B=H6<BdV;WNK796,E1:1==e#\@.;(GKARCcb3F[+^=G_68J^&b<2N(bJL=]f]850
// 2bNc,Xe(G;;YM_7W0=NCV+c/KfcQD,]+::RQX.ORF/a-D^4e??2^OMHQS<57>F6K
// 3T\#-#H31:d0SIg(A0(-Ja@HYDf_<-_6:_7/+@M[N&CFCb(W_&gJfc_[)+Xg6/W<
// ^N?GI@M,d)(c<)-((3H60209FE^b8CI<bT)7T=)KIO63X>cEG0NQ?2_>HXMe2MH(
// HD8aO?gbaEbY5KN,+Q_R]GDE2^AYSLCLcTDDW.5N]4DXW.-F2D\N-8;GcMP>+UFL
// Z[gDg;@cVR;FBVeQGR743W9\BC@G95RE?PfPBTaUB>B1<Z6Q3PB))e@e3MFS[ff2
// 9SZgJDP)2017Z?.:Lb)ef^bNbN4Q56>]Xc&NK>&fXT/:J;2-;>4\UCNbUVQVALQ4
// .,=UfI:]V@2>;2a51))Ea[O)F;4GfaL8H[-V\Ef7](,/3[#TeM_@KPQ88-<53USD
// S#;dgZLWPgPRYa4+cDdDF9SWS74g^E&3\)>D7^ffG=OO2A[7Z71\TLfeLW@3TaA,
// (K@#)UDN?+>b4X#:.1WHF\bJdJdd)JORKAJ/8\Q;HAb=C-CBRW?9#eL+2+J8T>(,
// d0-8ZUJ0gMI:-;X/AN7/=EWRTYXeWd+b>g&3bUa-(#O#Z^g#G5:-d02O74UKJ?;Z
// bX-(F^<e-d)08F9dS7TVOb??CT<[b(DGF0)6@\ODRb\]R]]?_@T>e3)7R>#68_K<
// 3bfbWf<IFd07CZ>)R4E9L_P7e9QXJAeUF#)#c^Pb76agG8,=;N3KRD@]^:X_,TFg
// GV/6dXYN\G<-Y.FYE5d6AQ2D.XYZJb(/dT)8,5OGCe>9T8M43EZfPT+@)5@1_#c4
// PcN@\),74Z^a@K<KKJH0?Wg=g4QeBSR^N#3A#RL@:[6R<2>fbL>/@8FT&?R2SETD
// 1)FVUGDEECFPMUP#_D\.b4R+U<:P,dbeNDSATdJ=gFEEF4&O9W]]=b7&,&2OLR)#
// O0C+gBD8UgLQ@2>6TZ.:b[_90-7JIcR26SX62//d:=58QBV&S3Z5T>Z>aPTUP]aX
// >be5,@-BNPH+Fa0]E3<OH?Md)@N\^KeT#+?9ZG&?&^(#X5O7\WB#d]/d:=7R<^0b
// #cOHeID&?49&GDa8/TdQBM^JA3IY^>)JgI_.,>#.+f=\f;7TKbc&JW]P_.GXE#dg
// ZV)KFA>]cI&CU(3J5Q/0+U]]:L+5e[Q57\@?UCRbZ:56b.&dAU\[I[IMU2EZ1ON^
// \fdW:,@F?7Kg0W.e[f2,Q\BYJ63R_7YfOYE6RW_VK5<EDX8UgAY2GbA:a<78g@O_
// +;f,,/)]952Lgg(41JgYO]=dFLL+Y9.SZ5OFF/THCDY81YRWNB\ZdIU_UaEWJ5?P
// WE9ad?VT5L5_.R)HEK]7T4UEZdY+g^O(;\N1D>(=VUb1MB,Q<4f.aK>RN4K6#13[
// W9ZL]8WKXO2X4(UQ7++K2.&@+0Vc@L+?-LRM^->].&\26:W#MM#J27)^T83,9bX7
// SU.@>/]+KeGH)#XV>e\XXQBV+5,C\+S8_S_+?:<UP=_@2P;g<RTW[f\?CQM9>bQ?
// 7_<0N87,-1b(Fg_Y(Yc/E?4OYFQG>&;F?<)f=bA630P=O[V4AN<8&ISNJ9=1ZMZ\
// +K]5KDf1R,41D;O]^E=e.FP(H+:4@ZS;KN/7]5]/>&^RD6.6XNOX>Fc/@eG-F6</
// <KW)1G++,PMdfF&e.(0&8d-KNWd,^g9=ff9JQ5WE5S?;(;WY3=>V5-H=Z6:9a(-H
// O>aB]C1]2J(7A:#.;W.AA,&Q@cI3f(0PWX.cC.:A),DEE5&+;8PJZL.b:YMcAgI&
// [/NW[_?(]B^CB3a;Z&K_671^gMW5&;Z/ANZ:1W>0M8CMB]b(_aAb3Z._Y5;KZV\-
// )-D]PX]H?4/]^P9YGH/C/E^>=W,0<PePQ3QV>J#eX/@PcDcAb4.?^MYX/[;<^/HJ
// 65fZ)MVDZeB@F86I]5X,-J7YZ2CV0Vf471:NW_AaTDE4H.(g2UPe8ZUJ@ZKXc406
// 2]#9P)O0IG)IOfO+fE:YQ4F9e)9A\2OO1,S)OA]-9EEd^G<^b;5Z4(4-\GP,E;MI
// 1E<;2Yc_Idd\T+A2\^CWQ(AB<GX0CN+#O:D5M?Z,fa+T&Ba:7>N,R58(-(#fUZCD
// QCM5>N>@&;+PLF?d1=,\Oe8ab1X[J[T28Z-546K7cG5GgdeD&J+Ig>X?9\N5Y@A?
// eU(IQGabOfcaI:]Y6[#e<2Z9?9]VJU9IH-9AOIMg/(MWI=5Q+Tb>]G-^:2\#)2O&
// 7GVaL/^Z#dI8-A(=V3^A),OD3_]_?KW<+.Jc:]B):E;-R0?9/O#8ODBgf(1V,cHO
// Xg#4F374)>RHL:H59a:JbJ7?W4fP,Y](Q(^(N,9(+#R?A08Uf1S?TJMg]YBEW]:;
// #g0ZaLCRS;FU#(33?;MNYH]32=K(c/K:-1e<E/0J#<F7d&M#Na=[RIaFA(=Je_;F
// dW<EKB;d(GK,O48TCdZ>ZEF//8gf^=954I40Lb32;W1GZGVgI-.V1>:/]DFbBE[H
// A@AFV8&Ad4H3CNL?DNMBFd.&K#&YT3V_e:QPBOOG/?F.C6#.9,-NeeCJHT:e;c<6
// 4dEH^CLG;:eXc<&,CXVdLYXeH]Z@A/426;d,YPL9cAg=5O1PFN(5P4I7E@O=Y\=7
// D4)a/c&FBMAFRW-U,:<0I8+A8dEc-),Y[&2[b)QM2Zbb\_M6eZ+U=e2K[Q(\T#1)
// f(_:8YH1d9SE+I<]K(Hf7PEgORB)>CUNX0Lc)NWc4=S6H,NN3J.g)]&G?8Ea:-FF
// 7&R&dFZMOT,?RbS2V;<0Q+)6ecY;6AV9?3G.^Pa4P)aKJBE_DEVT..CPM7]K#8=+
// d63g;1UVR9Y&X-&8=RR[5AW\+0F0DY;<eA9(PNAYeESBg6B-;K\NWBKgY_;[f:;&
// Z9P3Pg,ZQI1e.Q]9X631+Q.K#]\QHE[HHV\(MgPV2aHB\f9_U]6/dQ3H&&Lb:^Mc
// 8^g9HeK<\0e-82H-c=c@#3J_O^CX(RNYL&E+La:gK9).;R^+d8FUC3\CS_Y4b@Bc
// 5:]-;2#L0LZ])cL5<,>e<c_O6C4,T;#<;fEX,8);()-aCY70Ud^6EB_BeY(?c0;W
// G^IO8e&)g_?X1c__eX,7KLHbU=G-UUJZd1+XU]\^a_W/RKS.A.aZP2LG4U77SK=F
// +:0U>WMVdY8(/MK)+>P;Z?4I+BN8eOX0=K1ReG>1<c.c1(Y@2aE6B-[XN+)@KH?4
// (#[N[9C@/5OA7-eQ_@&L.J43O[O:(3QR1M^:GXB)5:5W4PacEF1dagL;fD4WT2+6
// ^b>;XB&,3:PJ72a<>Wa(bID;R3(RG\f:?@R+N:8;Xaa[?1S,LeBWPXM68_U_dJ\3
// 1C6ELPg&cQR6YHfFL+B_#S<:PSAP2a&_=4;>^95b15,@2g>e<fP\)E2PI@8<5X.0
// [f8(a8[,:_FBK<1<H>e95-B4-S6S?448^+5YN1Mb]QSUCO2cZX3X>+(\5Zag?5G<
// d;^A1QT@4e)T_8/)+?S<=KC_4)9fc/SBO)7[2FXb^L&Y9F9TUWHfXJ^fF5/a2bCZ
// C42Mgg5)ZOaag#D0)9)INN)K^L,909HDc?TXd<I8P8/aDU;,#>b3VR0gS87N2cKW
// MZ0L1gX\_.eQ=)CHGPea3>U[,TcHE84;<Q)6#L0;90@eQ/3bMI,N6gd.M/QBX^/Z
// 2)4#@K]FN)+2JXfZU^g@De5MaASZTb2H9OX#OWf@YbZ?T]W7.@40;_[?M1GccY-=
// I0;8gCS326Ja1?:DNJ/4d?GEO+_)DDgT:9Ub3PW=/RHYJfa13?[-H/4B=E:Jb]2H
// 0SE1@,5bG:d&>GIVJ:0G])QO5)\_0Y:3.QOL,0K3cW?2)A96RP:JD_[^cT25B.I?
// HL4N<c#(4beN/,I44=ZRYIYJUADI]KF4U.QR;HJ:9NMeRf3?/,CaV[FN/dMT>C<W
// 5(3P[Y)K\g+<N]9<:WN_#TMP-XVYT1<\N,;P:QTUd,MV_&[DH7;NWT^#dL(3+Xe0
// 3[>,ccO2D41g[TT_(9P.ZfeM2\\H&?be=80]WFLWUCHN8ZgE6Kd;VM3H9D(d.ZK;
// 8d\..(+G5C5>EU\ae:M<1,4D[A8+6DHYe->(K0U7A27gT0A:\c(I\4GR>O.)35EL
// [D-R^/[a.))X4?GY1OLLUP(#F,TEPffJQXW6CQg+_N+E18,2OOUI3U##dZEW0HQP
// Z,/D;&+eB;Qc7Yee2bbU@:TT_<N=/BV1:.g(\B/[#gAF<;fUeb\XVbX/6V4/P)0,
// 26C1,8e2R[cPXa_KgHeS.)AF,aP6X0;TYe\WaN9;I>a\QJDQF89fJRYPCIf#R]+)
// TJ5E&/CU_Ie[E4M4EY,2B#CL.83JMBB:?(:H4A]g;<D>Z,d,Z)Mc+]2U^LD0M3/S
// B8+_,fPB(WQGcWV2dPaL<;=&19.XJB?/[:]aa.<S2&FdQICPUc_2FS@I?O7]->E.
// \S4C8-H3@b#d;>F(]-d)\[cbFCME9^@,DM+FY.337G+<IO/?>:4N4I675<=6?:IH
// ^ORMJbF^I0KVReba;;dUC>8/]N[7X=)I+CA/A&]4e&C=e1^7^-35AJP9W=1S.TT\
// bcf2]D<eJ83&-1]g62J<b6H=I:X<<\(D,QC(@S.#1>a)?E1Zg,A#3f;0eUTD:cd_
// JNO<_F>9P]fRM8^A5KaARZ3:BI^dZV5(E0aSY<;g]c9&BK4YQX^FLL<FZS,FH0[K
// 47)Mg9<YC8:e6T,_dK0[K4WA0Je4XePaDT7PLF<W:]Dd/:1aT[6-_^RMg>HVgJK(
// EYYdFd.]aV^NCF8]4HAe?=WB]8.]]=D6IXI&;b3CB=fXJXb(W0dU:^K60IG+LQ2H
// ?X5G?M(.bV&:a;?;=0Pe/S<1D#>4CcC<JJE2J[MA0-3CFT^Id1R8+<Q[=A9XE?-#
// (\_@[AL,MT8eH6-fS1P_\7G+#8QC>->Q\>>GN/[+@_IfM[?T^27Ye>,D;)c4H>RA
// 1?C5\Y>EHWH=KIB4(bg9K0KMQb?;;5ARBN7YAJQJ#dEQfZ:K:V(I.JG(SH?,HK)Z
// M4QH9M+c6S6MAY#CgI[G(>CG(W[3;E7W(PUcbU_O+;e8<ROa3KA(W<B6B_F)\VCI
// Y]g1]ObfB/X)O\g_#V^YG(Pe?C,a0_/Ug2c7B[[5<_>DG0^a8W:RX_62DW:aK34^
// FR9(d_F3-3A7UZHFS5R0Y=]F7,KTJ]_?b>(S]7Q;3JZ[5CSCfK:aYY4G_G3Lc.Pb
// S=C?,IHAXJEBdS0UI)#;;87CB6Hd55Od;[,SSGUX@3/X@?NbGKX[W1U2d3a.?Cg-
// BLC:K/_gUd-RU;+K/T[G0U[5T8&[?B9UL_FJ8#9f5c0:gHXJ,gB6/4Kc][F:9K/_
// ?HR4\Z^2UJSfcF?+U?&;@Y_c_Bb=/.:-;RGK?.GD&#.g5.SI--0#HP/K7+QYF]YQ
// Y^_HZJR6BZ@UD18/#7X7QE5D94WLY)?7,V,1?V=Q.V1bH1GIC+YbZ(.(UGOV8d@X
// UE)=:T8a\3:>UbYe>]O;gX4\93XC#LN2C_WDO1\DX+8O3^eA?3<U0D/^b=\=J2-)
// LWHWV/,fS5]AS[dWc62]3_bTHZ,7>HB=K0?Z<?3^-4?P)W.e,OIfV[7g_&\[W9>F
// F8_YY\^QD\VUVU#@#TcVK60>#2Z6)Db0N96c:.GdKH,7(CS#34VZa+QBMgMHQH2g
// 2<7UdR#Y@KER-]I/20VAg-^NXB?73(KfV1)49<AWBLT@JZ<A7Na[1P#0\03PdMV8
// P.1)(N3XSe8773e&AMSSMG0SaJ[807?Tb1e]P+]V>(9bSH[gD=J=\fQ_8E)R<7(P
// WM6]b<KDI@65YZLDYTZNOVFP.\4TEDE(?8M<XP0+0TVc4N8:J/CB]E#V;c9]YC7)
// Sf+cFP2EX3];9NY&(65F2/>9??[+/P<O+[,bf+/QT)E:J+_eb&QH)Z&W7-G6ePFY
// J^<?Q__TQ&&N4;(6f6:HL?bQ\3aa3g1[V>:/:5?3WWO[N&PeFW^?U0WH+Dgfg)/e
// L-_?3GbL-0BQA(;,SJDDT^;HK:,c_Y^.]4;7^2<OG7#N2XJaOAN1]YgGG8+eK&DB
// FJ#,4&GT,]QQeTS&FHMO^1Y8M+O#J9]Z2:#Z-V3+-N9TU?@Af:2DVC^-BO2Jg[@1
// BQ3K.]e:_MfRP[[_fN+P^Z016Q(@_V=E+U@PKVSNH.83@JfaO=gbWMeTD-FJN-a=
// 9,b7HY,\VJ[:I)Q0PHCE\X46\,JAB4?<S0+O+)bKB#S#INOE0<c+?UZ&9?7e4f<d
// -NCM&9K?7/2N3MN5CAZISB;/e>Tg)?fL:Y4-2B\a5E^Z;&GBMEDZ-U:(<@Z6G=a[
// :ST][K0(9(X0C4[MB?2E/:fVKWC\#OUXc_;WdW\;]5:/VeTC@6Le_g[8dI/c<T6A
// FL(Kd7Fcc4LDEP#:TC_(JB&cSAA@5TR\:(BCf?YWC9&b>7]?5P0.8WYZ=JJ7.5E=
// =@HaD-PG-(d:\2\VH[@_Ze0._B7O1OWF1gW1VKaN(+C3TOE^c9LUdXPeA0]D8MDB
// N?P2AJHTX0La8G)]G&KZ/f6SO&e&D.T=+N;aP3;<UAH^e;/b?Ad>U/eXL)/@5SG\
// 0FMaV8ZJ&JbWEMG)DT#a3]]1d\OOF-,.[;F)Wg5(;2,#>\[\+&1#@0)g>SOQZ+XS
// T-07S3>d(W&Y5dS4>cA2f8a/\H(LVNYNHYP^6T9c@(BX6cXdDGWf]::R<Ac:J?-H
// F_gB9a<XIK=[UQD((d.1A9Z_[I6=U(9L>cgDP,GWPJ//,2#5:7\P2@&HDP5^4GLT
// &:_-b)g++d2^Aa<[?PF^XM2:3V7>^cAD>UPP3/eOUgJ.PTAb]7V(NTH[?46_)/N+
// 8(bGH:H9]N+5G-gc;1H8G3FadGM=I?g.M^@N79_[M(;(a:73&S:]@ba]aL_f\05e
// 4gYIFQ\Zfg4)S=aJBf#=g3H6c5GgBV5B4.+Ede450+1YOXF7HgY=+4.g1^;]7;&=
// <BGCWHCM29,N4S4aOLXOYcYg&Tf1M=\#0YQC)N\(8M;A2KX2;OcFFc<&JI^I)_19
// RN3(:B?NI+-?+&_6#[2(SD92P8BNKHSR8O&TCgb>gWGDa#\AQ7D/M3W4#)]>W3,A
// 7D\--7fg4\[KIG#D7e9g^e[d_bX<&ACPP:_/E+C;>)#2OOaS@)F:5)-/1UN;b-5L
// (G447<4;73=b?4=O42YN?O+OS^?XA\QL&Gb/X7^(,GLMKVCS9^=5U9-M:M8-R(K8
// @b_ZC4gC[KZ-G7GfZ/8+TcN61f>285de)2/SHVFFg0Z?_Bb;V=]aIWLVfeF(90.#
// +/b=R7_dE3VOU_@c-Md5:Z+RTL:CZg9F7<>@?@U6BRZ_bGUWc+ga+S[+.8Z(+WaI
// c:a)Bee^,4]N^gD]dRdb,\;_;I9X.?_YTaD^WXYZgbGHV[/OO801;/5[c_8<2__K
// QK@PT8/YfSJT&J+I3cY.VC\?1___^,7JX2TgG_(49Q;#_75Ve5AOPP&f;BUVgH9J
// G4]T0EAO4c5[3W@c(@M/a0V6-(D[Y294(4_COf[+La^7_6A>)?Mc=3,E6;J[.;NY
// X(VZ)SB3BUe<M0_;58\K<5g-1UGI+BG5TKCPb#RX:3;/aM8@:(S@#J5D&:W?S?)d
// P=T)W)6&^.Od,F<;_B9E8@6CW.A9?N.Lb/VF3N+5HE@])@gJg@d=?OYE4_C:RHHG
// \DK3O#FG\U;d\ALcC:8B?\T,]e^-P\,^5)0K:F/JIPWbca@L1RTH>g_=c\ZQUF_4
// 2P=gDaKW.;_9OaBV.2OdY<(Z\80FKX?4/46L(bHBS(c\&fT0]d]6]^,Cd;?c(5G9
// &W&\V;Y-^&SJZC.UQHM7A3#Y;]9@.[:=#^beb]A4;FNc,>9I^PgWL_.ZXWU:f9.2
// Y:+FKHa=V_f=L9a[CaW9a=]W[NL8F#W&\(46Yb<JYeE:C_fZ)aE=WPHH(^;W8a[J
// [8O>H]28Eg5-BYM^OYKZ/c1;#-6Y\@+60cS41P[WZ4(;GI=:BR(D+IX5]4J13TZ1
// V[JUAKQ:(SNe[/Y2LEPD?Z5[.;.fa_.?aH7fYM9RM,EKD^PZV0_ZZ)+P3+:(/?9=
// 5\OL7_879R3KeZ;dQ;1=G>TA^:/?Gae-VDcd-S&;ONXJaT->-\],6>:^;>?g)O\=
// BWHa]T?0/OP0#830ZLK.Sd/6G3B,T6F\V=a4AY/Y9d,d\WZ1P3&Q,IZBfWH_dfK_
// bX6?;:Pb>=+2C?(=KK7=HKA9Z@XC_A.I7GLZU7McT3IgQ4aU1UE-U0\,4a/E0EDK
// :GD+UTWY^4Oe9?PVf#9N.F)c1#XaW_BbcSNA3&f8XP2S&X.TbSDDG[S&b&,_C)E9
// Pc_(dMfT3f2=DfF332AS@146GSVPM8+)XYfa27&SKM[f-4&ARHX/K?2_XKgKPP_^
// bC7D0TN9g>GF^g/fMd+ZfR^9+S9.(V=WQAbE1c+/I=@5(bc/#eT?BX#C4DJ>eM2S
// 1N)79<AQcLB.]V+GVdDTYY+gUG73YcCdIP@d6^C[8EW]bL]1I73b.L54fGB-UFP?
// -05^Y)4W^+&EdSCFTGO36?b4LaMc4dEMU@=.=VVJ1BCKNa0(8:;JTL++XGL5M8g>
// a,bA-H/e5@7&,1G(NE3>7:Hb70@Q1g=S&>e2fE55+4-:_<g[^&52PK_J0WD2EX_T
// O3aSbR)Rc?@CFVD3BKH_-B.VO8WWZ^4?U5[DQQA,?^G(\>aQg1HOY4RWDNe\K;Fg
// ce6,PV&\K:ab58eACc1FMVXOa;:gJf<2g#H<SS^WIW3>PO?^RTf:?VEdR.e?L2Y+
// PS\2;S,9BTSFV1)F=JXLN_T-L=5HN?b>?Y2dS6ZH]39A;c@2AbKI<3M_BaER5]Y=
// J)8^?NJJ]PPFFZO5URa[ZG:<T)9[AG(J..YY-WJc#\1PA8/E&=a+@1]d]NP/2=,W
// dSMe(Nc;),g,GXT>8cQb(.g5A9EG6;^6ZNDLS;HY1)KPdbTS@:8#94-8-\7#J9I>
// VH?1)_U>\P6V6M-U;:96:TG>>>+)QNZF3&#(V>HeP2KeX>8NYGE(#e\WW3TJ#E:S
// CN01ADg&>B[:/=.WEDZ5\]IIc.3T>H1<caCJBF?3c.-0,HC]?+Y()TERMa;,Vg(L
// 9+VOVX@?<2T9PCK+E:-GE@fRO\VU&#0gNZG_5L&egbO-Ge[RB<019+GCFP9ER&2(
// WOX7C<\NH5=DGM1A(DYR/Xe.;,ZQ&c\EULNd6SS0?eRbWRY7a=GE-(TQGB#L:a=_
// B]&F(?46N/Q20[(b9SKCK,=+.2X2&K<SIM],IQ#=/;PUTdV63(Y9L;3e/_2cR37b
// bL,#^N)K)aJ>/5a?YK7WE46L3]/GH(BZ)8f(^PAFUR7/6ddGFJKfd.L7\QK^BK;[
// UIX+27S3fLY:>g7HUbXP\5<[TaI42BY6#,7LO@]/&XW^Sa8R9JQ3_TSOXK^X:YU5
// bDRcGDO.J1Q3FF4d1GO/<?,6E2fX\Eg>TJ1(gOI];X&,YTE:>J&OMHC+FT_^aHS=
// RAB5<IeDOO/PR)fTZ+2#B3DeeI#bd_gK7QC;YUNV,<Pd(dXD3B>3WH&T4c86IZ.\
// PIf=af^CQT#0S#?.4<=C\U@:_3baLU]:ZdCTa#B;L@)P]Z50(e,ef?8OOB>aBgd]
// O-R=U<Tc9Q<=#61DJc(ZDeR:f(XJ5;Q;8.JF6OM^U+f01RX&YWLg8O^=eS,aLb?c
// Q_2fX-X.\3?g#]B6e20bdJYR_f(+dV6(4gEM^G;?-3Pa8OZ]^+.^)3DIPJDO\7RD
// ZWLW<P.T;7_cDWEeVgLEG>)B_KYe90V]CIgM2\LM_,=#?Q>^(Hf.:g^YF2U0)d,V
// ZU[@S[_NgN).4=:?:+?f]LLR?=?#?8;5YR0MAZ6GWP5aeL=7a;Y:T<,7?Z\J9NXc
// .AFT?]F<ZE7\[^H5F(+Y=_N+bS&@6[T:EZ&:0(5Ude-R-0fB:.[Y_[YTGb8c.MG?
// )=:aA+OY9R61^VYV=U-SI^:.=K>9<UMOO:=RA/7W6G:[YUGKC<M[Le><<49._\FT
// T(N@Ib0R=07)6&6J(OEI-^dJ)[B&L/JB@1>_]cCa7fdJV5LDVP;390d1a2WYM#T^
// ,H\;Q?5[6gC.gVT?E6SH.Vg_883G_#/ab3g59c0fQ+/CJ@Ha3R[(#f=<7bMMKEY_
// RF2_N1-b^=bN;+80P[KK\X+V(EBP;TI/B0SBGFU-P9&X;XZ+_51WIR?CO^V<U19<
// M&RH?@/6#f6Ra8QfV/&@]O-QEOb<97\=ZcSY]a6<:53JG<?A@=9B66T4D?8K&bJY
// 2]UYK8&JV:_&fTMZT9Rc?N/>O-TOO1PM2R#?NAZNIfCg4\[WD=4gRQ(X:gY#IC:K
// ?)DP>U+0K34GF7TBS/CVT)-=3I[<\I3AEU)(26[E_e4P8g2cQKZ?Q&)H/LS2LaMN
// 5fHK.H1?Y>Y<IC/5=VQ-K3F:[HM>3(]Xf+.D7+1W_@8e^6[R1Q+I^/6a1=7ZO_)2
// :L5H8UF=]W2X_YVJ?a\Ze8LO8ACfQe=69_BNYFMEHAERPS;?OML.^+O\T80A^2Y[
// MIBdbWaY:[NVF+[((Mg8\PEM6gDg)5FCWJ[N>)K_SR&ZaUgU/BH045&B<f=D]=6d
// >YIe/USUDYd28Y]GDKTeD)c7dEg(dZM(=Tf_B#>LI/(DW<4G&M6eRf9L.\-dN-O#
// 6=97B6?JL<Y4CLW.G4U@6H\@&9P.Z1@(:)K-B^/(1AI?Y2?O=U;7Ee1GJ-PERFY]
// :2c^2::PGA5fbK^O2842G0?#HfX-J,f>c9U<OfRR1c,:Y)ZU15KQa1_UD5;V3IWb
// g^NR^&+&9?271:@6UT2:O55FYCZSY@4TPH/A4W;&:GdG/99X-Q]5;:F5I>[bBTCG
// FUOUGQSN3e5#@Z2QS3aO;#4Q43.cL^,;.6U5-1=FXPfHG\/4ZS8;bZK)?9;N;a1[
// 0.eeDO&(7F05c-J^WO74CRE&2]cD<<F&S^_6VPL05^ENGTXX7EeU&-1;a&Y,X,X?
// 8P=F]7VQE9MMNW)D[D9SG;Lbf);KA\<3EXTF(3WG_W?,MN((.+cB88.]5fb,7\V_
// A4MRVS190/&aa@G&ZQ83]4BF]dYO\1HAOHE[V-II28A0:C:B[FH385C8,aKIG+IV
// B4NPM0@\+b2gZRVYG#ULPU3X,a3fI:SW6Y_;\L#2TU-4.\1&>,)0E06T.?1<RaQ,
// ,D8E@g<Y=MRS<3,G3U[T_QBg-9f?,<#Q#:T_>;FX-+4=.6HXRDR;T#IU/K+d03HP
// _L7.)04-b^M7M0cJb0Sc:[^L];,229(\98f:6Afa&ZfPNgHb.I-cD=3eH@Z>a9E_
// =HCa(.YTQGG^W[,7]4-RKNL=OZH8C\H6C@OOZX<X[5?K-Z?+T_cMWMB#;/e<67=Q
// 2WXIDG](&)0,CZAE3cc#+ZWagJZ2fOSA>J/6f@d:#7/Z\MDAZegRYDGR8CJV>gR\
// ]Y>,]:8@9+Q7O?AUd?/S+N&Q_4(8McRFBCaG/\CcRR2X[^d9V&][[0DE_T)AW;BC
// )E])BG4Ld0c9fU]DP^Ucd^.a:A[?a><G;CZA((Eg0=SINLX@&C(aRbI)aAeEeUbf
// @+AT6S[f0>O,ee/V<ZUS3TMY/C_Q_C<H/QV8@9B#(_2V<YW\VP+-DcUU,.^Jg(aO
// )U:#gLg_9EXZ^RXeP:fLJNXB0-WP-^2c93AQPJeR\KVL<[e]LggK>B5-MZ3D8efE
// IHd@e5/aL/H+d0T=>PZJZ+[+N8@RC(#7?I6LK4_AK?cZS-\F;;A/6,aC/-[c&?N.
// ?@aC;B73f.a:+9V81aUg\#S1]9c73AMT?82.@F764348XV4S^=596<=d\^M3Xbbg
// [^Y3Q?5+<;QZ=#dN-F0]XM\.@KI5;05_H#JN2LWL+XQS51f#G;DO_<.4W;<23K?2
// D^M/SWZ0[9#_gdH28KHD@2YIRH(21PZ?Ed+K(<\E.eP:9BG]8_T[)5cF_1NgKF;I
// 4V)E-.aEDM:AA1>XFY9GDPIPb<N\D^9N.e<<MG_5]aIAP@]?UOOWLc;1F\7(gW.c
// 3[:IfD6-DK0>3^VJY19>(C:]a4;?/aVCHWERO3G2G55MO4af\O]4>NN&9#0RF+3S
// <96BU/RgI2;7OIFVK#+CD:8(XQH>f4P/D^RI]LZ+c=>R7H;Q_J.<(KVKVPN&,ARF
// dF:3g&bdE7U98MR@e,_fFE6HG@[M@)0/6]CdANd.Y^\.f^M#[;G>7#f?7X62D3@B
// Z,8=I0(D=:EDG1W[4Ua-<Z[+^>X@=PAAaRKXMSgEY>g_P2,?_I&HC.>XfJY\\c^5
// ,RCLRM9OV<9DX@?D9NY(F8bHV24J[?(^T<(M)WD_U8T(.RPTIZd&=e9=P@.W[L&V
// 4c?T30H?Md4&&93UIM26E:(aLN]2.WSZQ@HG+H6O[1/-:;,/+.AcbSJ0X)U;b&Oc
// >Y[gc]dBOJRZ.UIT1/.GM#-P6ZWBcBAfX\>K8=f6QH:6W=GIQ?Nd7F5KPO[(2W\(
// 5EfGaf4e1Cb5F[+&V>/^?4FDN6PK&8g:?&C(M/XOEZ)8-]SZ02c)1Qb.GM^JP6=c
// U.XMf^VBgR:IOFBP.gX>0RJ5@JO@,T&NPcTT1b6EC45E)96f;#X8:CI,DY61G&G#
// 9U#YB7Y<Y+bW8?MADR0M3CdYHZ,g[32Y+EYT\TM:S,@W]d=U=U,B^M/#\C;W3HW1
// ?a,aFC(\/U:8XO=F,[aI5P3^K]).001^a/?A=^LfR^R+cf6+.KKS::@UKbIdJ_R?
// 7:,?3>eB4a/^/8+4d+E>N+[?>6I)fXK_[Y15G:@X6SH<NB7)NE-BM9TB/,O0=8>U
// [fOR<J](8^[fWCJ7eKS>Z0MG50)e,E0P7(SD,(fQfT;g,;86&g15K]a#eDH\[)IK
// Q?HIgXgN24e^9PM,Dd<PbbN?.fa+2TB3ABT3V6IED\e&NA><e5R&@R(D>TF\@B+4
// 7S^D_M:>=Xeg?bREI1;SJDEACMO2NH-C.&:UF5QfB09F83_4\C6S+-/a7+AL8:;f
// g&.S):[)Z<\b.HDBFY6R9-DU-XQ7CcI8?QOX5S0ER@@RVZ#S8L??C/34S?L+^5gN
// 7#<[,cF)47OISa5Y5I9J3a;K^.)gVA0SLYYZ<ALE2TU),LZ]4YJ>/aXe4LF@D2[E
// MA5dg)G0-UO5IAGZW9a60UOI-,YQG7^:43O+SM,V,8C1.VfWRIT08&Va;9/@AGY^
// :&^M/:<c__e/Q<)[[IZ?Me]O#[D&2J0KB^[-A:Z>29SPHU(,6)GaIa/MNe)RDM?/
// O02SQ6-[<,?)EY7A-_9@9e=;C.4We5B<WEgL:6XMV[0f7aXG6cH,D5Q5LgX63UfV
// E))MFGfW.T@VP<XeF81RPf)[.BN4f1b+J)8Y&_eSM>MZ2?7\W4C)53U@=2:#7X/U
// &gX(JOKUC7VQ+[^<,MOHDU1&c+A&cfK:Z6G#:C(0Z@U&fYK9KHW+?IMWP&B7?(9A
// SA(KF.?bPW2W(eSc?X8EG:+Y<4F[)TRNb;\b9D0CQZG;.W1=(B#7-<SIKCD:]gG&
// &4(8;X0A7PCM40cE>e\MS?bQfKJa15YI8]M>8=-5cP893(QAB6)?W5V-f35VIJT.
// NY=e^d(d<e:H;80bHa\\&)[]>c-eN__b4(Ne?X@P,AKa+8Q#Mcadba[fNX)GXD;M
// (9a7-D8:FeKDU4E:,@<UddX5f5]a.ga:Q+2QHg-=9V1V)=@P8_+f#FG-<1+S0f0/
// ?^25OYS_4(BNg<K6.7?AbKM//N,c5E35JWM.?G)PZW4\U#<EHA1D693TG]UQeUBN
// 1JKF;=^NHA>+TgI=(9K8;.3d(0L#H.8=?7.PM\Lf0Z^b@Y<Ba:1Xgd>C4P(56R=<
// VeL@b)(Z1I&AK[]P&4gbK8K,b.,U&SO/>Uee0P#1&S];QH+X:ZecG2^:EUNT>XFF
// J-;>NLc&X6gBPIZUXGfNACAIW\1=Mf(PB0f0WC\RTN/a\0RRNISIY0<_QZ;(D50Q
// >f:3:b:<RIa7_PJ3RFc4=1Q99[RQPRIOI^R\\,c=1\.e_6]8&V>\CCO6^>173Pb;
// 8?B)G&\13O,U.]7[@,U:Yg\09]96<8)^L:F?FDMKC@GQ(QL7XP-_V(-N0+Ag&UcX
// f;CT]7egJ1]^+_S_T>/0].XDb\ZED.9+OA.F4DSXX:OHI(1[V/1]9IU2(VLJ(AQ9
// O.ZA(daP\X:W2I/Y&;Xe&:&5GGTVL1,:5F&(&XW]3Hfa990gd_7Xf+0D@Z4:<UA7
// ._d1N#_E2-.YFU6109N=bJf(d7-:_1:F-D7_)FM[6VB<5AV(D(]I#O>I0]7(I/PN
// F:[7)#08YR2;U\MCb5R3X9dcbN)e29/c+2.P[Od4/RSXP+QJ6)4H0H5UM#W\(54;
// ag9:1)LR/A@_@,H\\;[E4I@_),OK,U+J,5.S\DLWHcHf9\YfW_WITca@Rb4>8/3K
// K\@:QFER_&JW]3eHD<>fH:64(<NH.ZT\adRE0,:-[edTZTB\2OeRCWW[,aQ-LWG^
// _0IC2/&Q:L2/_]ScX3>(9I?,FeB[[WIQLPS-[V-ND[S9=RCWRH9R&Zg,\.M)e6/.
// BZ&7SaMb?.=QB?9,&#9[c8D/N-,E.KOXA8RWMG[Yg(^dR0LM1\?A41ee]L]#DVg6
// D1<PYccS__+^&Vgc;\VA+?a,#B=aV=-f?IK<W_A#S4VZ0+5Y9^#M7d@]O0FB2BaM
// FeKc]?1NW<Y,cDSc+G-Jgd2\2#4Q,F8@,I5L7F=_C,M>-R_D_CN-4&.Q>8)H-?,5
// F]K3<CS1W2U=0R1&_1V+f,[LDO4f98(/4_E0edGT^_#2S<9YeH+9W5=CWCJ=c7Ad
// >FDBRI/F-G\RbQR40X_QF#TFCG@>[TQ;;=^J\d=82:JE^T>bMJN2@>Yf0>A?R@LR
// V1\&W>K=e6RDZ>-+]1&)dSAUIEB6\(]d?4KPbL<W(\L&&8G9AbGB_60;JPG?Q=(>
// 2f018?F;J[9^1_JU?C6V3=ST8K)5aN.cg3P2f,5B/@A6]:/O&5_JC4F1S^aReV9=
// \Z261JQ=3S&ObP:3\0G?4:cE8^cV-OBB_@\=G6\@I\gA+W^:f>;Zc.H/QTfY&a2/
// b2+X7LZc(-&]b-Z.)3e2,IBP,6;GNY4C;gOV;Y#W>1M#K5@VIYg^(NRHbB/S0--O
// 5HFLa#R4Kb]._<e^/^Z6?Xe(e&P82gP;,9c][UDS1TcBc?+:J4<Q51.gcfNPEBME
// FOH/Ec1))RW1>5&:7<47[@O1K4YF]/0gB4GTcL_-4^?;^V)Zc<9ZJ&VgH)9.c51)
// ecDNa.3[1@EB9DVQXAU.aL0;HO0\4NL;N;HJ[RT)A69U:[]>4\CaeP:9_Z,[6aC@
// TQ5^[.PaF(B^S8Q.Q1:e262M6QSSG8L-=[6JI6UT_@=/Z\JUN,Q#_-WQQ(L>4HG=
// <9(B(2cb(YVI7Y9#N,3A.-1J;.^R-KCA.)B&2\Z::cCV,WIF<]F_K]EWY&)<X(9Y
// .0I5f:8+[1=D3b^9\<TE?ZZc;[HRWd9f,V@f2?N<c]eO207IIW))I3+T<db:L48N
// #3EEC@BVG5b<Q,3SZ_D[2e.Y[GLDOWAd)T:)#VK1BC5I(f;3I,=-+6;Z79_D:0?-
// <<&/ML6PHb47L204F-d1ZgAAPf>e54-2>SR0Q-3N-3(S=8C3bC-[KZCM5ER,9\/S
// 1)<Q?+Xa>[(SOWFK;HcEf,g8<4P:0dH(aNT]:U.2<ZBE(QSKN&YNMXGT>\WBVcg)
// .bU\RS78d#d6g_7CM(c];cSVRf2A=dfRQT>Gd@;b#g-GIYb5]6JQ6YC3>/X&g_9+
// VaGF5c#bGQ4\P&cI=>?-;Q.4HS@D;7<O&XVDEXRS>[?1#E4;:0>+T9dW:6\OW[[;
// 1US_cffZF9:4KJH>MRKT24?Ua)+EXg>J[B]cgJ1[ZC^8..G5]Kde==XOJ@9I7d8X
// EUTXLFO\8J:>Nd&7((P@TJQS5Z9WdGAMC=bd=IdW^.b[M+6aXWHJ<Z/Kc2WY)=7/
// \74fUYYCeH-L<G7Ke,B-8+&0NBFO39fK=dMR^)^&GVWA(0QV@7(3e\dX\g^0KFGW
// ^&BR+,27#5Z(P)3A4\YQ,Q(#8]afGTTY@/B+aDKO@(BN0V^O;IA[7B_D60Q(9e=W
// c)6S?eVR?P5<16-G;\ZS_fBe/,\S=Y8T8>_3^^OQ;WcVS8MK;<VHc&.S\9083;EM
// >I[;@Q5+<T-JY]9R?8=6;E=+;:_.fgL#(74=W]9aB3&X7)A+dWHC7:f4gd&+(9C(
// :9aAGcD_O#.>9_Cd^C\6;]@K6BdF?DU]]J;Sg[A[A3PJY7K47VZQ9/QNW9Rd/^9?
// dgB)2(75I3gI8=5XQG-8ec][#:6Q@]H\cRLVV:QQK+Ve(dLV+6Y.[f)33Zf[=\+D
// P+HbZN)(@Z7FYIfO+,:H\TPWG_8=S#\I5@#HaVL+4g>D1d)<5c7?VKG_A0=>gN4I
// X;A^MR)Y,RFe/LNZe#C/8g]/[LfK7(CHBD1DcLQb0A,L3Sd^-QZ\M^9OS6FT@7YL
// ^[Y&:WXWf):NMT<CKXQUKVTKVDMF30PS>];S&K2F,LHQ5]R:HX9QGQJ,<95-Jefa
// e-3W?V.U//HIW&80ARR57Ncc8#?RP&Zc(UEDaeO(,.?g0+Q^9VOL37HfV;Bdd3WT
// ),#,F=M5W\<9KKff:H,)<Z&D@C@M_8QRQ&\C2HQgG#c&YEbN;.1efVY+a<&#1DMV
// eEeF1IcgF&4FK2DdMFY=g,1R)f7LN0IOBRZAAg#-&S;K6XB-07d6J=(A8XcJFDNR
// E=PBS]RVY@8@g\5bQ+1N[@]6C/N=1Q_,b/A<5a&/(P6JBCKNUK,ec,Z=f2Q;K>W5
// FTLX<gS=C8eQYCVEb.XdTD4Y>c<T-S[9M,M037?(&PZ-RYMM\3S0N.HeT\[c[-&W
// MY/B/aQCcZ[McC?>?9P#TMHRL\DeK88c@8OgU?DK4&WY\HU8;DZ)bQeL45>;W/-2
// /a<Dc,,b0G6S3^4\a.,\5T?cSKe[0;P@52cY7J8PS@0<YW)]W1/\X;g8)_/5:)5?
// U_C1H]^26;)A7)+W3Ie@AEdH/^VS)E^M(IN,>&:SUc\.RC[[fWW3=b=,Ngd;5]EK
// eFP7:X83ERPbV(gK==,.T9EGNAG@>.,E8;,KW6SIH[W9.g1G?Zf,bH<YV7\[F/_d
// EUCGacV<EOQ,QX-+^b@AMY/C9O>^2>OUT)_[Q\]LXEJ&+4b5R\E;eZ;-HFH;WPd5
// 9.X?ZGD@(\H;++@67GB;<)Zf]UID.gZ+B[?M3e0XMIUF;PKJTM4Gg@V=-==&#4JD
// OCBa<b].O<8[d&M-C02PI_KL]gP>/#WXF>;GUPRc;EfA:</5.E^6W&_8CV(LICMF
// Z_Qb7,P-^gg)2@M,K7HA9?c^<\8A-5Sc_,1:C78_ID<1;CL9L4Ue&Z2TS5E\Z-<?
// SbX?>IBR7?GBb@[e0Dd<03N&>0:V/Bb-8PM@:f9UN&[OFZ;ZJ4VU\+0S3/C&8\ML
// <#YY-&\0Sf=8S2PQcE[dccaaI49e79aMV2;8Z:TZ\=Xa13CL]F0]1#K0U?_SG>G1
// JU/82]Jc:&5c8RF7^,OBJ9I],JZT@g&fBb<.WXF>+6KJgIGd(QJ#0NN;fZf@.=R-
// &#fUUb<g@L8]Q_,2bgFNJ-4#GJ#HUJ13<aB@WfdK^9XR4\4-29WNF0b.,V?c\RPT
// 2YFa<Y,;a@cJ3Q9(V^]8eMC@I?:J=G]aUOW;</=SLeQ1K.S6?^QM)f](.WS@;Yd#
// 0&^d@c=#)2gSc+[GHU2=\\=.R_E,(NNQ/WYK04G;&&PC[ec^_493>R+g@R&cR5cg
// Q0GH[&f8Q7,@bRD,&VgVOD&+M^EXNG0?-#c-RXB?f\@]\U)(cNcB&6R0TM^=T7QT
// 7(TIY3#O._3H44WZf<9)_bKT.fZg@4VL4P/1N_A4)]MZJI/PEM@5F@FZ_\Q=]5c6
// ;H9NT+_/L9EbY]B,,1O47;DeL7cC3:>PGMY@L3^FF5f;GOZOI@10)N5=Ag?BL(S7
// OTT^e^+C1]cD]Q\L0X/.:2HX\&LeQfI1cg;I=8&M]R:F<F7F.LK6E1<8YMZ?cBOZ
// 2#_@HF-A1S(;9@IJ.;_d+_DYP6Q^e45Icf8d(Q4+@Nc;Ec2&&);IM1g]K>[7E4T0
// 4-(LRYEK=69DIH6L64L/-SBX:EL01&)6bdB,;GCI,F;H_,cZ=YE1d?V_7DRC8Bd4
// SBU?,)aSX??IOLKd=5)Va8XA3ZO/\=>VC?C/XZDeX8gSC2.>2Q6bg(_VN&_JYN>1
// ]dE>J-BX\IBT#c3AK9I7?cD5G)@R=@4@7T:66F>2/-T4;Z+I);#SBE.7-+=I_(N:
// d;cD[6NQ6V298[\34YYG?I&aA[C3c^c8E64LaZ3G,LN1[EBY2HS;F>aS]4YFJE7G
// FEafL=<S#//c>1Y+X>1BF,-4#M&Y,;(@B9;^G@J://0WP[5\gU-.8bMD2#D8V06R
// RI]@YJ24)KZ@.YagL1,JO9(R5G:/QTc&f2#P#(K58>ZPR6YDATc>E@W3T4=DBNT2
// (:cGLe37,EQ&1.?(9O4BQ9W7^b9A8OIJfL+?NfVJ@_W]e4_B1)),4dMK9=QLTG\:
// UYI(SOUJ>PS-Y,2C:g7e91;cV3:12(?[C55I0E3NUGVc:_<Y</?NT7?g@+&,Ia37
// ([^5<+;81KLW96HTUKY(8+9&#.(NRe2+V9eBX30][7Z]2\DgcX50S)9g<Q(.Gg\;
// EY3\;AS;d[LSdLRN8N&\I_+Pf0^BbR^]ZSS[DK@TPK:MNP_,-f5F0WG6H&9QTd90
// FU+(M/30C:/1Da;T=aEB\J,/YcH4.\gL);T)01)#e=./=FFR+^G;B:,TDD0E.gVb
// 7?:&4d97WLKN:NC#+=2^<E,HF&bgcYZC^=gc:OZ0^RPO_P37FH3O.cNQOgdHO?5[
// _57@Bd@3U>YeQ>9C[a8=Q:FKfIHO]Z-Ig:-1()/c91(=6JIIE,U/0VS33,8FCb:@
// (0[(J-/gaI.d\J=GTKCc+HT&00g3E?c83ObLB&4bWfc)(ZgM,(]H+C\._BGJNRaN
// 06RU:.H-E9A5\;f^8FP6H\.XfLFIRT-[X8TPE:_HVbIRV<I3?MG_>S;_1JLQ?L];
// &9\&/C,Pd)C&fTLD/FHHc5EcB@+&391c45eXVSNX7Y>G4252Q&8KG):3JebXM:@G
// b(:M:F30X0V]&TX-]eb:.U8[ETbL;bSg?dK/\UFf4DZR79#fU/21[>NUTX0AI?KT
// 4.IeC_E,>7#^JFHUF4KN+=A=;:<f;X#0b]a__N=+WXW[C;OX7EPHC)QbbEZU^Wf0
// =fPaF@;0EM?JI8Gdg?_6[+g8O;U,b_>VSWL\efe@?,<Xa8+378TdIO#8AO(f946a
// \RXaZRY?62a(F4W@3bF#f]dZ(=DWO;DTFC=gB]U1XUEW#?+4>e:/4]F4+]Y]T038
// ?MEEE[Gd(N,>X91TKY7V37g?7M_W5(0_-[dZFRgb/.[THF#a1L#(]Jf/;T0BAKQ]
// >(F2_f&?M(579WAV?QAAK7VBH49#)W227+=<.KS4DcP.-H(]fSV0ZF@@]<4M\g8M
// 7ZUgfd=U/1]P\+M1C.KYECBd42VG@1[Y\OCa1FFb,<VgA@&,aa-dWcYJVRM.TH#R
// @G^57_.D8dX^JJ=(NM/2ebW7?Lb^/dBEW7)M4ZZ?IX-W:XOW)H?aN0(GWQf(GfWf
// KPfN?A,]:ad4dgP/cCHWf=,@&RKQIOKcA6/[+1b1M;:URNOgb^_M2Fb<@ENWV<.4
// =gMZ>J,^Y^GUP-8)X(WJ??M[0?dDNC8M6D6=dXgIbU]>=[8O#fV;<RYeU(S\IS_W
// C1Z#4Y;#5^]gUURC2f(G-3-c03,GTTYW.#7,:ZMYWQG=&.Y=EC1,5HaF[Z^gNCS1
// P.9E@.V3?LdT?VC><O_5L^>TBB,RPdSAg,+72?/?V+_\-?EICW4HIR4d-G:;JXTK
// (VV36[<M/KXgKXZ22a4VTXFc&aZY=fHH]T3IV^YK@a+7.5REPA,79^_a4):D?DE9
// _0&>_+WS?<&?Jec]XIIUe8/8[,<9+#,N151?ScgWIL+4CQMZQ>)g\B-RUOX7C#@<
// e39-B.B/3UZ2/KNBIFUWK9T<U6[aV2V=>V[^UM&XTQcYIB<1[-[(S]=8);V5[YR-
// &^ffa9>Z0,Tc\d97T9GBd?e_Z2<D/Bg(9#XS)(8-D)fHX->LaKJLeQVPUXH;e;.1
// ]=NFQ3DGERAeE^),I&fP;\b)A[(>+5BB;<9]+</&961L<)WS\^#,A00cUOW6N#0M
// CR+#-;FT3G;OL])>J61D&5=M935AHN_V.1CVYJHRZW/WFf[?c\+.LNV?,4EQ-,GR
// 3E(/68@WeW63ga.BK38.Q]Z;Q]>)S>(BY#@e[A>G<SC:bB_?/S4?e?9g4;e.Y@e1
// ]RS)(H6.GTe8\8f,4UUSDO1@M5^;?M(#bELZYVG<-a;OLM<,SH^0&-YF;?946A5X
// 5[]L5[G#S<C+#YHFVX&#>]+W(V;XBO29N:51G38=\9-<X;=N:a^>@.SHa^WAZ//=
// [\\TCM_D^](dc_dT<2:[TFGMUd=dY&O#,[U#=I1M,5)a?M(=G4J0gVH.7/?f(_:\
// UAdA&^#B,8\c.ADCSMO^@)TZW-WYVGC)\-R\g)C/,K@=aG6ZY,G;2MP((4b>=MCV
// (F#DGNUcd00G3&5<(2>ZNd0\LSZFFZV-c5]W?-@HP,VQ8_RWbW<9c>2:]Wa8c3>K
// -g&1bXg+JA>)d?RfHUX5[e+[-4W+Q3>+dYVP6YQHY@96Q>^:aR+I.=NeO7f>:#4Y
// UYGAC-Ve34H/>#A.2LK0>ML;O>38:\AGT;ZA4YfL^W+cRDED6Mb4EQOX85(g@c6C
// #Ug[fbJ[1(D4(].\^U#B]JgINT=<\GB7Qc\[aDV:-51L;gg034e(cI.2dg_(KV41
// AD-YOfbbbFcP>g\\)V:J6&Ma@=Y#=ADZ:=fU5.aP,M^JO;/ZRW=NHUA-7:_X\V&X
// 9AA5H1]A8_<TW9BE@P6[;eA[N]E=\Ea(CY_^<SJ_^V:>,#Hf)3(a/Q3?:I_6^+@a
// ZP<YY/a-<]YOfN>0MQ&5^<U&+V.,FRIQL-SDYe;1E.6SLa13;cN:?dXZ,dRXBdTc
// D_HE6KI^>@B3C)/E<:Tb3<O\<]N)4d\?<ANV4g3G<(DFD)fKAJ)4gTc+4LOCF7Z;
// DTb_<;fM3dD,Z@YIH01IK1DDM6>]A,;J+b]1PK;NFV#bAD:W0cU8OcTL2PT6+JP5
// ZNZB\UXX294Pa1PZ9Nc2M2H98Yb,<4dc[P.fXe_XZE1Z0LHG^74[]LP[2OVc2O3E
// bOeO;^RN5N>eDe8^6X@g626NEg,;]4E+,S=cP^P6NCMD16gC5U#&Q]dda>G<S&8d
// UL>-9+8Je&&?DbX&_RGP[2c8@N/CLNMN>LO)6WAVF)OgO)7gb+8JD-Yde7<0Uf/H
// @^^8>gNa>LVIVWc4\\,bFd:BTIb2U7.HVBUH66cZ>cRNO:d4E?>6<X0(.U?4CC(/
// @M@T2BaN<N\GVOGP07/XHE;/-LC4bb:d35266[B<c;IOBT&QV6ZECgO0E;/D4]1P
// V;A[5;N7-DBSC]/6N62A.g.HPU\ZMaCIF3TF&RW@Z/96;SD]>=-6-dA(+P-X]gW#
// ^0\Q>d1+3JPS-8gS0#NAB=D<Ze_QOSHSgA9JVOORZ<dN20Ja&K,RBLV[VTB4WR0X
// &SD0B=fZAY^\8,2.=S+5a8.4F#N7S5M#Q2d)DCF)Faf7,=E&Xf7:N3=[eJ9:SO,X
// >-^J<RN+9@I#fJ-\W>>JMa&OM#5TF3_TQ\EOOg.MB0J?O1>c.JFEQ>:XY+fB<gQ[
// 3233Xg;E\,@BZW:U:Y4[Ye5N4BF1Ge,Z#P<WXC#[-]FS>/,/<E5E?X/1#KT3bDG;
// X-gPdB@O,?eA/L@<7#,&_Be?5..2F5baB&ge5K]e-N8FXSNWE@4F5b=15b3NWHe(
// W2X(-A-gZ(AK6Z&)&bF<]V;=#BAQ?Z^O_/0D/+L&7F2HHJ_MI(K1IN.@(-7F=Se@
// INWZG?KX/S?#QfV8(\_@9^D)/+JR-d/T17O4Y8g6\2g+AE3@+e;aW_UU9]_L:MMU
// ?NSE3S(3e]75e&89F)P-=#[Vc4#T)C3\#+HA=Oc6aJ<Tc_cRLPTaQ,S]@Jd8,U/a
// LG8Sf29H]<b48[CO:Q,.2X+PANXg[V6YXL22_7]>_^B8WA^Vg.(_@[eN-dTWI+DS
// eOcLFMcHR;@6=Uc[T.)0b]I-DR-OH:AVK,:TP52R=&##+/f1cM11NXI,0=SC=A7P
// 3,UA&^ZTVA+A)H8;(9\H[Z+dRD.@-[38RT0SMA#8gDeOV;AXU<XMVM[\4OX\@48^
// gfGK/>.UZH@QH_@<_IO\Fc8/d3<3QHH0^#S:ERNI8XJ-X4e1.A+,QQCQL@\8^<PT
// C@P-3=,\==AR(5CCVQdMH1_RY47G84VKRLUG0:I.XTD/8>L-b^1g#5N8TeC_OJM]
// 2X_1FA3dP-8,(YZ+9XS02>0&.7TJA8KSK+fVECNe>Y0L2UN)?/;e&RP\R;6SN5)W
// d5=AA06f&N0&PA5VW2WE9-F-TX=]H3O\ZMOOc;N:VKTZgPBR^4JDLJ[AMV#eBWf_
// E1T,8V&Q\CJW)PBEW=)=#ae<I<5F&LcFOB49gaXdeL9P34WN:A9Xc)P/J4H:^+EK
// JR0<N58HdI:0d6G)9.]8=9S_-T<:FQb768^#Y0Z#_^O/@[g;R1BH:0\-dbdGec\=
// JRIQ[Kf(VA-JL_[1P1MXB;M8cTC+3RfA-?&Nb<\N2bHT7,4M+F]C>R/a_O+US-)f
// 9d)&:K=083B2FT4H0XI(5Q/Qc6MG+#V5QU9))Z41dW7SXecLe>ATEUOPQ+5<MF3.
// [S.9PTKS2MXFG<?:W@0Nf8M9T[K7<C<Z^[\N87f><g-_?.X(8[U/\]\a#??=P?<-
// 6H=79S@9)BWKC.17.ScC<eIU;.XYbaWCI&&O]B.5YN=4@6O6-./X.F<@T58[7LQ#
// @):>4a0YPYB&[X<R&9+d]7ba4><54#5PfB>K[L<OA0C8<e]NW(9gY@#WWE(,?.?3
// bQTSJ0]=eZ#UH+X?)]_H7cNDV57A1&Q]?Dg=A1(D8gG4;KJ8EXT7M^WgLX9-4D@^
// dQE[10<O@^/,VS(a912;a(&CW\RZ0?a-2[(E(b1C?))1Y=a3TO>YL9:V?^cYaTS9
// 7g+HD3OEa\Pd17d/4__AAT<a)Q-HcPNd57Z8aQ/XIfab;XIIaPO(MKCBAX)711dQ
// 9/W+8.CQ4=A\9K5c&:U+>/KW@_SPN[eN70PY,^5QSOB:#N156L_5^6/K5Kd5Va^/
// 3PBTGRCbBXEX]d[Q&4@2;N;gIQGOY+0[V@^GT96ZM)QTBGO/FD)g8,HX^=P\W-<U
// UFKYIV(O9?1H&+GK9Y,53/\S4:=52S-d#Z&^U2YM&ZO?\[O&G/R.gG\)BHO4gBU^
// ;=g,29HTD0&=dA86I05AY0X)J:]dUOXF]090FOT^&I[U5<V2F>EJ#E#d48[T+6Ga
// ;LH9IE,).+eI(XF&>PA(O0fPP-SdV<-D@Hbf:gG\f<e&^^FKNdNWJ6Yd6PBE3^MA
// FP-[AAW1Ofg6I^W.f^UC6>(]7QPGO50Y#?8?(e,^-V382Z&Y00VR3QLHLcEg89NV
// 1d2MV:fUBe,_&&9EfPCRS<67X>GV6UR82TYG_,^G]@a,RZEE>QLS-&R\cgc]DBa>
// :Wf-\+\8X[HLb^aS?TTCI-Q-(E^4Mf4UegY]a[E8VG_)R[J-a<C@#Y:;YFRT8\QL
// g>eG/L7:ENc;O=Q.c08DJ24]=6d;D9HVC2cX4I]6Db_J5P9\[?[geQV_TIf0eD=S
// +WKND:#OSUI75#Z-B/He7L99G^4S5f=bdZMS?cS(KY&/KZ9.WdUEb50MBeLRaRF;
// ./e[,MQQ+N=A+c\=.+67MLD/#N:)?S\\VN9W)W>2B)166-E&2e,R/Yc8_g72(TcH
// WVW6?URJHfEU^=fZD@2Jf^41Hb-PYJbW\+2Z.H^V^J#Y3SegN+LB1[<eH[dcT5#,
// =KQQ)24-Z.[&&)9]N6b>B.M7gUP2gY,6dA1:>Z88-+M1Y\R?dSVW4\](J8>IWAN-
// DRNa?(:H8Id0:.B9dMW)W=RYVLYTO\7B/1&bCUZ6=.Q>>U-#e/HQKg<C/.UD]H0,
// c@Qcd8dU04W;4M2EL>+c-E6e[SF4A4cO+1=cc.f[=XAP8QPbR)[ePeU6dN3.LQe6
// BJ(b@b&-g[Z@EF[O.H]+UPcC,O;B@+Z,O]GVUS3;-bR25TK6@Q9+?05Lf^Kde/eA
// UZQQ7_Y,IS2\X/8MNO.8c93]Of7Qa=cG7D@@-FNWYH^6\PKa2T1bB\(#Q=NNJQ@.
// RIZgO^117@OKee5I@g-4SKF3WJ_-Ce6.#gG3^8BVE/C[.EB0M2R#Sa/W)RER<9Zc
// EX3S#?0b,+-a(WZ68VGX@+4/-SJGAb7d=?SFN^F>;d#B,\A&RC\P<DW[^F2/B>.V
// ):\4,LPd4F,_\a9E^WHVBV8BEXg:XNGI(GN0O1>Tg?4e[5:2>X\d@U3L6,B(KM)W
// 8fa60=G\,@)O,N4DIP>M>S=V7K&E#5<b-.F.Beg;eWN?T7-NP8##5Me_Ibb6(Mg[
// ^gcUP0<F;-FIH7^N&N?R1KUT)Wd1R;D03+9STU6UFf_Ha-9;<C8#+\YK&PN,UK9D
// F/YbPOJ/>/7UY6&AAT>30,Nf_gV,Uc?_38?6>8DOWcJ,8HL_X(Cb3M5:Gg):g_3M
// 9V0(>QCaCYH0a:X9DLI6JC_M(QH2XMg5(>E\b,4VU@G^<#Q\P7&C8I?f1;.GVWEK
// ,e36#R\;P+]c8TXfd)@d-LJ-?5+0KSX6U8H-aEC,(L>36]TL_[5QbJ7g<#gI,33S
// M8#>[R^HHL-3IG-Z)Y[d+,/E:f0K^2fOAR=dQZ4G=A+^6QFZ7H?6:7[+Q3_-/6J<
// =52AJ9[A8-CWKWJ+@3>7:@X-]?bB4DBWP)U1;T[VNV>3OL=;bB@]>KADYL0G,LK+
// g\3&KdLK#4[4YX(RK4_&d@F[.H9T=U:BR4O9O3H#eKD,YIT#KFF#-&;_#T,C@Z2M
// -,94f@Sd:Aeg_CDE?a6/?&QA/C\N]6YBLcd0#M@0L_LYcaNcV&c-^Y>3>>SC)c>-
// -;C9+<.5fIPc)24#==-c.FRJZ/[a<#=bN6VfTBL5L--U1G#3XVBb:;Y92a_NYI4L
// >&03H2BU&&_>3ea1S&654.NILFU=C,>P_U)EK(>4dXgA=CA6>Ya?I6VD6^LNY/3>
// YU;AG3K@U4fB1BPOU;+_L(L?PQ7<.6NI:RB0Rfe5>T53XKDDaX?[(.CD-e5RDGH?
// E/@@A0L<#Q52b\9eZEH+X37bTNZ4[eLVVV3B<Z1a9+gEE8f)1ACWD.+D3]\T/EbQ
// =]U28:@1ZW<^GUG3fWX_-1+<.,RN7-B\JgL?,H^bC7-,/2NCAUgY8U38-::<JYFX
// :,1<-?@BI</G^T7U>N(U5,#UHff:];.0J)^#5=W4OgeGARZYJ^XF#>SC<3fD[9MK
// R)CP^&U>^[c]:\:/&+fJ&bPO><E#&6:X/UH7J;]&1dD0QF;V7_(OM0bXWK,@K<+b
// _EL2eW6agLW(W^=X1<geG&@&Y.>&Z-bXOTJW-Z_Sd<]6J8ZX\WR8D=J-Y0gcY-E2
// ]gg??QR@Q[XJ:GB1:Y;^/cgRc2gH@6>B#=6@]eaGBE)>T4U<gYXE0_FO3Ac9Y+^@
// )1M:ENR]QTDI1SV/PAU]SJ.[W>6.DEe;a>QVc4OKEfW/M<]DKDSLfZg.fRJFb((3
// OZEXU]YBS<e)@?-7:X#=ZROM&I+;N[S^,;GF^,:O69W=eK:g[ceL[-gLTaP1eB_.
// ?<O>=SId14Z/SGgJ/1Vd:CHEQ\#G.N@7XU=K[fJdCP47gRJIN7F&FKf6\HU^,e8(
// TL86/c-=2YT]Cc>4R>_6Y3:8dZKf.-=0aeb2?C>KIOUM[d:Ad?ZWDW?;JdbebI5O
// Tf45MK]TdeKAF;P-E?Lda,(HV9A6&O4&UU<EegD5+3NQ+\&UG=56f_;_.M=;O1<e
// gfd)M(E[)=5/SVQ#5HO<YITD;R(R(/3B^PN:Cc\O_Z75[T\AYM,<]EZS5UG>88V]
// .O;-JAFU^Pa?J5&SU?HWN##gU9YL1Da>0]6D<OS5)MBIfU?^]+21;REMgeG&WbP9
// 6fTDe?2ZZ#D^&2cfgZ7TIcN7;P4^WRS)H@O5eG<D>d84FKP3c816^\+W-^)E]>RO
// ?4RM:DVaf@HRHfWSVfgPE,eVfNP;,:fAGW?FG/#SD9\B/E+:1TWA\3Q06SITIHQA
// 2?7Gc\BZ;P=@Q>AV2;UdX,5Y+#[e3[V29C78M^M3REg2#N4Z#Cd_#S/2<@YI,aa,
// L9?FKN=8LC\Z^UB7-8F3Q1QCL0JT8DN6/SWTb_G.JfNNKM0@&OX/LOI8Pe[;I[G,
// 0#Qc#gUU<d4S>:Z,_V@-Sde0@eIK.[&\Rff]\6PK?)Fb)G,WYD]SCg@D3_cAM&8X
// \_G_D8DMT_Q[[DH^-D5-+<Aa3G^DM\^GO6f47gB\VX\/(3JV,)]Te,PH8dQQ2IfP
// RXXU6ZI_WceC4/YJ;WfB-HR8_67/H;,=C30AX@1Xd_IZH#+5[KO2W]&SWG)?(OOX
// OYe6>R_cU@I6P^>.XX1]Y&CYOFLKQ^^+0_#WRgIW60/=Ya:J.S?76;\DU40>cL0B
// U-a_>ET7(g@E3?eTUU3NG[/T,E=:CBa]F/&J7bg2@8;a\19JGO4E?B;JaPUB8Xf7
// Af7--,5PcX05\DG(cA2(]R8:K^4TLR]cYAS_RD8<dN8=+@WOg2J/ca)f:;H?):90
// 9]MNaAQ9.:WYAgZG]/-+:-?=]ddgM4S7eUL4KK>?Z==(-XB8f;\,F>H;G8bMHQf]
// DV4OO+1MX1dVDJ8E<:06=-53S1VaD;3;T72+D;Vdf.e@V@.W>eAK+Q((#OU^g:Vg
// bUQP;QE1B1U=].SDK:6D@96F]Ug2+U:gB2\EdIeGgbGA-]E14]Q-KNK.fA#9]9D4
// VYa@Ta&/?e(Q<VcZ<U,?7e]92Z0#d0f9a#7W)^>FPYI0)C72Q=FW=_L/H3C\^F&6
// EMWU\6a:eYLVAGFa#I4&&.LY_5e+fP=1Z@5MeVa^ETFL5:4]U>^\65Ub]RP,9N(Q
// 6?UX?F18R796CgNZ7\Z;2<5:JO]=@GG48J+S?@)1DM@.5TEAN;:RQJ</bJA>CNeg
// @bEW,UVB^SVXe<LC.8MJAY_YQB(\4PMf5XNfFFDV?F=WY.VKC&YbYD2)@VY2f8L3
// Q062Lb\-^;T7K]3&7-Z_fK27RY=I)(K[/S5)]f.QK#ZTOXY.;=<PIC2.I:#Q&7XU
// Z_@:KK^d(5,<g2f^T1K</<?&f)<LBX/,OGH-9U/N;C+#CN[RW9AC:K(,g0J;GRSA
// eg4)=;O8NU/_8FS&XB]ICZ[&C(3/Y/P6Vb^Z7E,a?5WE>B4d:H^fT:^<EE&Q(\3&
// c[^JKT/^JObNCa#PQB(-Zc5>5?]G#g&AE-,US8fd,c80U461dcQgfT>-8R]/&/>b
// +P]/^@a<;\/IAbB>ATY4M:>AQ,45F=KJ?ZA\-C3e,5TS6S?AeA0#Agf1g)[=UGSd
// 6Ef,DFW_Ida1F4g]BONR31OU8,QRcf4RN&<e/1=O7.f0_=g_&6AgKMZ#&MaHDc[2
// 1),?/:9FdbVcLg9[_(&\Ie,_L0-DbYYfN16b0JZ#0f>,?[WOG.0gfBY1aJNWKdVe
// T3&;9c2=X:X43FDF,^\HZVdG<Y7IB5K60\[Ge<VRGTK1;^+M)K3-?eaEG/F+CEc6
// D<0=)4B,OP&NJ@PI9<CQ7=R=#_.T.g?GW=a&[Y2Ye/DUVL\eE5=Y?D14fg6FaVbG
// S3G5T._Kf<R;7Y#Z=T^+-]+CS?;OL:Q9dD]P&Y22IQLK4L\Udg1(J.VBXHIQbJUE
// gIY6A.>.eT7IdNGUVLc58WEGdJbB,[U?DLP0.RT2(R\J)\e4KCT[7R721fH):74b
// +]g+[-4SCPG7/U/E=cT+[Tge^TB4Zbf?3N[VC:ICG.B:DI_PJOZJ:3IZ4)TTVdV@
// ?+#+,XPVJ[g:FB,L)b<QUN--YcK2fC06TU4ZEFJR?MONCKHKI)P:bZ?M#3O=A36Z
// 2A#01<d/PIPXQ8RA/OI_\G=Ce=V/5][Xd>,5B,>L;XWb-D3<5:\46(SY5[&VLBQ7
// <gY-/O2A.ZV]LQZ_K#H8<KRgB4=D9MPY1>PJ?E28]QYZaPZ,@0C4;LgXTTCgIOH&
// 3VEN;c<R]_1@eJU+.+f[6,KGLH2Xf/AOaX,e2/?0dT=),f[85TDFHe.F-^),;3-L
// >:;NZ4EZ3Z5.O?N.BD[4eOeNgTLcGWQ4\3f]UZ#@d:(\8\-/YK76LZPUfXM9KOCe
// JC_;_+;@/Cb6X^JMVbP_;C]);XDeJY=>Y7&99/#gJOE^CHM8.)Q:7\GZ[#K6\\PV
// )@B.];_7,g_\59b:+8/5YON:4M^bGNF[5Ud(f1U-^+W;@CU<6Wb9Zgeb12]07+=B
// :X-Y_RD&YL/9M[a]XJ2FH<^c,KL-OC37g]2]e=4/Oc5NJA6_P]+M1C4S2IL.QPcZ
// OZR149<(@_[RTK(V(XY;9g<WbF)YU&&)Y[.XTOW<<S.ZWEebIe^#eb(@7XNMG5[]
// g8Ee/2N<A80f@/\4C<f?#;YVeY0/MM6f:La:RAN9HaE1aH-Afg>D?W01+^/Cb^)a
// FdIKcJ,&8fQc)a+9F4[/2,,GMY.?_>N1B=9SfPY8_U[bP=ag/T=<1VaEO@GZ;=FC
// b&L9<&(KXLHP@IG-Na#@JfJW^Jg_CT&,MUgP4@Ec&S=H5,2b67MO6cdU^(2[+URJ
// SI[aKZ=KDPZUMe9>Z&\H#2O^J?NO:2+NGR<I6_e@L4#OKT2/Xf=MdMX1Yc+4XBD7
// a<Dec2?9OFRdG7.UC,V.8KHLJ3a+b?;OKEb]A-)H^NWb(,CMeENF15_S=a(1A(-&
// SRKIN6X7TFf\9PIOT8()(=)990MaZ&4V7@a]+DW<cDK2f@DZ+f,ga<\V3J_4I:8G
// f3K;CK+-#<X:T;?9-_,.\eC\^2#f,]CW\94,YR6&LS@T-WR5)X]ZOQAV@67F[LE(
// PH[XTN?_2#ZPd[Cg.Q><aGYb\LbbS#Q[#;;U70,,.R\)b/#cF[HE#AH[AN@OHLW2
// W7]=A58O)G?9F599WAC?ZNP]BE#NIO=_g^J7S9^HB&\]#>S[^7/]AH9&A0OB-b^.
// +dC<#_aVdc6[<.U^Ma7.d6/S;]J9ffcJDAL;2775A-_CJ:E(9.UPcR+;1E\3J8^7
// D/#-)fIM>)=ND&5JOZPJ1RV1b[)6>KVH]K[\G(c#[^C?Fe60DNaD66)-,I(dIX>I
// 3@L&]>g9O_Ed73g,;ZUHUDD>6(B^4QZRUT3-JKN]g]X^T4(RZUG\^>.QH<_XeCM2
// ?HSTL^;&0\FBVOTCB^3RIJO-[@LW(B7^+VN=C>#>g:(bcJX;@T.IQ9f#8>99f+YI
// :=E(2Ba:0<()_8aWf>^#[(dLXfI;d[S2-LeP)O,dR\a+TF@BQ>K9411QCZWZR<8D
// ZNBX0W#SELJBgfS?@6F@3@)e9=gcQ-PHSX(@B]BZ7D4^ROX(O-L.eO/]@#H7[_KU
// F;;0ABf.(a3OLG5-/G[XHgfLD\7&gYJGWQF;GeBg0S@:QRU=7FCg,;<_NZefH5c/
// ^LRb[CW56+G(C4DL-)OE<DP95eQ]BMF06@^G>LYWK/1LG_HZH/>QT/.;#YfGeX,G
// >]X:/K1/5e>&-VH9O<?GW##,UKY^=HcY5a6)4WCGR8.KX;#^;;@HB8P3b[4RRQF7
// Q(3bcH-Z96>N>265PO8V)OL5JX4+^#,K3@Yb(2/g4Jb/E1g8RQQRJ7F\2;)LC;-<
// ]?J^-0ae-fSRF]2R97)XgB]172\(EJEb47J0Z[<A213>B.U6C\PZ1^I(U]3<\0HA
// ecP192?c3W(Na3c&C5Y0D.gD0:DBLJ>N)TeA@dg3\??#_^cPN9.P(-/)85?H#O)E
// aE9K[+W0.LWH(.-GZfLH7c6S+(J)4V?.LcCTg(P7.504gE>=MPA:<PaNNd2MX3XA
// .Y@N9)6PK7EGTa)+a9,b0&3#]c@a\TOg9C^^Y-TMJU-aa(L+8TI_J6ag:1=&]GB:
// &<2XIZM\]2WF7?dU+1-A6.T\89;OISRY+-K6MBPH<?]<N=eW?6aKM=DX^gP9YOSS
// _?bDdVPK/5bK^g&e;WFR_GI:V^QGM3?TPO1:/gD&J]O/TTZ@C2<_DZC>PB04G=.I
// g?.UeA3SF]^d5#J8e4USPN]HI?Y,7P=/]eX7;]21/M;@cLU?D-E2,S@;^DfVZ&1K
// _CS,[K&U2@IJJLKDYKd95@9F855(e2JLU7WFR,aA7FBU1(C8:X:bM;^HXN@aK4ag
// b30G(@]7<.c57L<&3YPUR4OYB=A19]HJBZED6H\R(MK<@MfF?JNC@)K)eBQ-7WN6
// _Q;BCRM:6]2=/g-H(>:QRKA&_B.b;(4XdO/?ZWB?4>WIcP=A6Z1H5V0>?ENCCTE]
// /&1Ig_4J7W0SHDK#1V^5Ngc)7c?V0\Z#5Q]bY\M>2>QPgfNRgE#4G=CER-e&-cL(
// 3)-e:d]/G(LMXfSVL:KT\#CTO8U]-K>7E//50Oc+4]M3^6f992:8B)N^9I(3D]+c
// OLSQCbBZRgWJ)HX7-,5>7>W[5D>3dYNKWY;V8TQ^6Dg8+H\#bb,MB)aHeU[^FdH2
// b4=++I\<QV2JRXZe@SNK[HI,;aH[-W+./SVb:d9-SdR@GaKXe/UeY/d/g3[fSS@.
// D?F;94e7IUI\IF1XU07fYgGCcT)<R\UO25483A;#LR?A3fZWN?:X=W7LQ:eNf^0G
// U&X\1?Q#26Y)Xg&B#eLX[.4Ab5FKPJ)1Ab93,3(/eS8A6&g+#bX&&K^T7eU#4=-T
// 0.>E2W[AD:T_Z54L^->7D7-?)3GUI6]E9@A,J.922K(?f+-SGG^AP7cA1Y[)(c<W
// ;+YdS@;aB^E3ST6X2J,068--7DBNH\L#?4@b2J.[Z_UT)5I@+5&=-QWH)SXT5S47
// #b.d?N\][9>L:YRQ\V3R_]S0&:B\J\S6M\>>54,K@/]X&XXT?Z9>BaODe4B@-a-D
// 6G/PPN<=c0];9f#]O<affY>-eKKC1Y4IKZ03-)4.B[R]]N]8^YbVP0/,)Decf^@#
// <P4Zf3ZbC74Qe43E&C8QS2PIU5IJE3\M>PIK3N#f0XZJfEdB5a3@6[8M<5^P)R#C
// ^5#,]D5]:WG?]L7(=X_Xb?<<SfgVSP6^,L@8ES705L^;&D@\3\/P?Z)>LJ&Rg7@G
// TA1EHZ4QUN1M+3C1F:QR(AK4ZEG\51#KD>;I>VRJ):B]VR&Vd#cSD4;R[BafI:[6
// ^ZJ2b#0^BD;:(9VWd-961Ng#gN@V4CJ&=cJNH83S2SO)b;&LVG#IAD#I/&;AH4d?
// MTbEQT2\M_=CD]e;B^IJD&eQeaM#;AEW[B.O+[B-SX8I/R_]D.L#.24=dGgSMeC;
// <<WK6HVQ5I6D&4N6B?:+.JdC:,J=0QfPeBfC2__(S+GJ4?f_dPC5/KI7gK#Q83@T
// 5BP^RDS<X4ba],9PZXcD_&J4.#KNW<(K<+3N)=K.2_4FW>SBUN8a?c>\/Z34OI34
// 7J[P\g<QDUWQ:6O<GVUY/RTMa6&?RL<P?If1FQR&RJK0Lc^+c]SU.7e?FQ4MV8aI
// ZJ+Q4_a50D+c>H,:(O31RX(D@@X(g8RU17)UE]CaXYCb8N\3f5Q=VaTO,P]\S96g
// Hde5UI:f?#0^=_.ZDBVcTMdT;##+=e6GJ8d8T#UV&Q^+[_>V:@3e;J;^WLS_9E02
// 7M+CC?T@A5?:B_gCV#dRMdLIZ)56UTc]M.1A<U);bNd.eO\H/gdJ7Zf.?(Z:2C\c
// PM[e96WbHZ>d[]##^,6RHY^,DZ27;&WR=9(/WZ1G5)6J+5<-Z^+[T(6H<:01_7dc
// S[J#eJ,D.&54/PFV.\J-CbI31N0g[T/Tg:?23OGabFRNe=23<VZQ[U+RbCRAGAdY
// Y+R5P?A0>4,@PF.>V[[gRR1A+J^C5_AT.bY<:\4cC.&5=HDe5AY94;#+OL6Z-?XX
// <,I8^L4+Q:QbTPLa4]HY^\?Z9Y@V[8AP;Hg&ZX95I#J12+KV(/K:[76YfHWLY_G]
// CFe.9E_YZ[H,d58CY,[F8dGCA3^?TeP6I[0]#RYSRbg;Q,6L>_Oeg:7+3cC@ICg+
// Sd]:f7WRbMSM399g31GS<NA//&V7<<.dgZDgZ3W+&QAZ9Q?LgNT^E,R77Z]XfE\K
// 0[46)9]W-?IM4#L[E62,82+g]<4[X;@[XND=_-+A7BA3+Nf<L=[[]d<A<R:ODQ[c
// KKZ9O:0G/O>SN[=IV_W]6H.K&:TX9=N[d]Af-D5>1-T1IK4b(8Jg]QK7<O5_II\Z
// (Ed_9I0?_)6X;3fG2P_^Y@X+6JZQSMa4:?dKab:KKHP(MXB7?;?B>QTecSQ,N)-T
// Tg-+76?B-(B,@Q3X#eI:Y445#cBIg<K4XYIIf<8.c[G@_C6N-=,:X8QGd8+d;-+K
// &I/2ESQ,0>Sg8G5<afR+A5bVFR(bJbd2LNgd0.)T45G#&(DI:L-V1L7MX;3B/da-
// -NU_A1e]aUe5G3UO3/GcZ6NZ;)_99eL;((Pf+I4S..#Kg)a,f@,ZaE4?TZ-TbN__
// 0X[>-+B:<0YEN&9F<&4+EXb6^=Q/T,?D<JaW0d@G\@7#f2Q1;/KYdTOMGCA+.&V/
// Y7RU_M-PUC0\::g4@3@H6&dG)+3;TN8R4,XMMa&P]UH+)HM#0XKE:Oc;0Nb.]GgJ
// @cKgGQ);ITQJAH6\]5(+1Q-@L4ZK@Y\J]gH:5L1>=(d5C_1D>(5MA?.MJS+Ta=ZP
// >XEaG><B_S8@/.P@P(K+e?XZJ_8]6B,)U^>fc6]5VQEfSG#^EUZ3\L:PJD.f#;G^
// .4+VOBfZ9Bg.c4GO_aB7T4)NU+N);+4<6.5db&S.3GYYB[KJ0WG+HbOG+[2:BO2.
// +aD[4.\RF_;O1b859Y2dFc<[^^6MWKPRgC\4U=RD6XVXXaY3T@EBMG-@fcDE=(+/
// IKTTe8O5#@XQ.WSUBU:eR(G3LRNU/fR_H5(]P=XSA2<AM0;ZcgXMOfd)Q>V55A1W
// 0KAF6<4dg7IbJ#F@R<Nc;-M)A_I_1aDA,5OUIWVE)\L^U.KWb?5#aa5bc,6O2P&\
// Q5_Y^P&H_/K/BVcNf42W#/Y29(Z<[=ACS[DWWC5T8>:_F)>gO^44O^,1VL4YB031
// UK3QJ]d+g7@Ub1J/D#(ZY3,g7/gbJb??F&Y8E(]]G/LIKKbH^7>QW:-Bg05[F2#G
// <-(7;WVL]K7L^CSI-GZO73M+&-L)cP0\bUN&ZCDBa02\8@:N@_4C@GB;.ZPJYPAf
// RMYNJS>GcB-6^]GWQ920<]U5_F@2G3Ld.6TQO^cMH-GVCK:ANfaJ8aR14\6U?WJa
// IIH/--]UF7LW?OWMW7]C0(R^SU:TL]aMCZ4K:K0(31QM_6Se/,9AM^S;M9SK:Hf,
// dN@GKK&V?Yf=Ab)MaV_<R)Hb;HE_\WVV+Fe613(/ZLTLSKU#9LAX[DJPF1RB#ab7
// 2B2]N[MH._fZ6<.>OD46(3:5:GC]GJ_Y@^R^[M(\UANMSB?NO4P^@02CV&Ed(S-A
// a[g.[3A9.Y8gF)+#07J=cI=^Vb,5bfKCfXS3:58J_V/)&<,[4\K9&0)0^](M=WFc
// ,D=U^JdVc<BLL&&X9^b)H,ZY27aF/3&#eU5bE>a]\#CWN0OT83H[HI_3-C&E9BPQ
// WX:2A=3?FUE]eY<TRE,<D(B(_<X(N9FNeC@a[RQ540A,fYH].9e=4CdER0US[BK5
// Me?3<?X/bCa[/bXU7P++aBMc=S.\3&2Qc=W/;WT=D_0c54U#5XQLQZ&34L2&4.9b
// +g/;RN7LEM8.0G&6LU,a\N-]G@)gX(HfRV#^628ZXY4g1a,W:LLD:0&;(;83SR_(
// aEf9:F&I1U75UA[f[:5SZD)2AICeS9<7fHD;KP=_@UMFaRPT:aeK<66Ig_37.>73
// ZS7@?b_9](OQ/W#BI6dF6\#0V.A:SQ9_XW@ZY,e,D?7YMdTXY@K;B^IKJ9.?.2?.
// B:U\2f3_Q+&?PI)<B+KfW0J+bP0dZ:<<@A;D(aG_5ZR;b,R\=4=_G>2[05#FHK5S
// 3,aIRbg&Fe?D<=B.6b,_[O]+Mg-8;ZC7LK(2566c#,1Z,GMS#D@B4ed:D/_E.aJ?
// 5U<3KQZIaIaN>LDbS915\]/ec/_[R=5E6gD&(e/G&2ZNcbMBKL@,/K^YX_YR65^Q
// cC>Sb(Bgffcd4#C?S?KVPZ+5JaQ<SP9AgON.39<#dAFM1S;BUK3fYTCZ6L(?--+D
// P.1BJgbFAGd#4@8cSNee(0NRR8O22&W91UOdTJ&QdW=d,))5:MOGP5HEOe>S./6X
// ,S,d?OfRL[L_NPFP;DY9&TfH.bDCEJPQH-_.NK(TeSY#6]N)@7F#,\S4IH4_^^R,
// /2\NPCEYNPYe+fHb^MW,5R2Zf3E-cOO;LX/3IW#FP3L(YZNT1IFD2GdbgQOa#\_T
// WS(F1b0ET]GU4f1)7CD6H@Z]D#^X/fTZ:Xc3bg:b:/T1CMe4AT2TINV@-/CMF,Kb
// TT(.M7dVaZNW4f/Q9PeNAG<+eaX:8]GY>/3(5#QeG&X&?>]\0H[7XZA?CH[bH=46
// ;eG0#Y3Y1g\O(^HMTOA3#//g(T#d\=I^<Q,dd;d0)D8>ZAdg&..[)N4/:]#d.__Q
// [+?#W1E#0M;ZP[c5(V3c&:_]W6g,SD@&:+A,#)JW2^9TCDCNBE&WDf6+FcQH6JVb
// :_F\64S\WS8/+9aI1^9U_VJ7\]D_JL.-.6HE.]b67MJ3VA4R3P6>M>]BYC+A,II8
// XT2=J9Z@5MAK=@3AR49U9XS1,&(;L_]LB+aS]<2QK/,NF2[KPSYYV>;BdZ?e[9,_
// GXJLR]Q2aPA/=3S18@Q>H7&NA[@,0(R>\PM71bMK3Pef2Y-@^8(UMfgcP@_74(\E
// 1;cKKB)N6Mb_M)AO/Z79f.J0SW2J0J=#e]+&Z,@bHBF08IPP#/Z(,eQB5;NP_bL)
// O4GDI/.(13_XB.I-][DS^]=U46KRL+_\J.B1.-G,Tb,07I\Ta@<)/gEZ]KCVU5E\
// ETgGM1C:;@/ePBa>3_]DJ>6F.b=XG2DZ:Y\L8KKf+N/8AGE\dO(UNMO^Q_J/64ca
// 0PgB.X-RIeJX-,Lb-7C7b\\?L:R.ANV.L7N)fK[:_c[DTH@@XL^aUYD9Fe\AB8Ld
// )#f@R.F]TC&4\TZ5=/I;>)/gOXaR^ReO(^a^H)HW1bf>@\U+N-ZTg>J6FfIBbU@2
// BYJLN^[GU2Y^.42,Y/D>:H=4\Q,(=J/9H;5((1.e_1C6^B@G;7dc:Z8/MW<Wb?SR
// /:F86M.6;Q=3X+g5,fI.9ge.-XD^4aA=.?2)EVc3d.GTT-=d(+1:d#;(fRK4<7K7
// Q=M+9ARNBR4^2dM90+aLU+?Z6,>R(VRLG=6G(I6B@4dRYJ;VBX0H>0YJ1T0a28YF
// B^gU(PF>G??7&9RY+/a/T/])STX+LeAZ3PS.>+6&O:\/15c3bFW;8GW,f1Ed<2^R
// _YF[\:&1/+g[VaQ]BD/#9C&6FC4SP&@a;>(X97[DH#cZC_QH\K#OJb80[@:;URZ,
// ^/K2bE-:\7S)=D>YF[84HTWG/)a:&[;;9I7fNKHGU8<\)GZB[^]2?8I5Q6)W\QD,
// S1N\K:c[0CL2_Qa<<ZTVR@865R6PK69@GU;D@O1BY/4K&^^O#O:eIge++:E4^H=:
// 9NdJZSXSUJUb++KG+YFa]GEQ&62/\.R0_,2_MR4TaU?4TJ2W.3WB+8B?C<_<ZA(I
// X^J4:M6-:J_V@PE_EM^S5\XTg>=&)9?@+Lf7734Rgge>d=3:bTY]fDcRHSZO&aSX
// -857NbK-#XDNE?[Q(CL,/bO^=AII=+Qge882HQA@#X6Qd:O-0Q,L8#NF3T42fUHG
// 9\SIR4+BM2\X9ca_?TF5,QV?FHcJA9+_S<],X>;MbZ:LX4:=.G]E+5R^3f^Fa]CO
// 0C@c0X=[95a-8D3M<C;63/SWD7S?S&.:caXEC-W9V#Md8FYTVN4,b^a;&YL.(fQ?
// dKdOb/;S@)S^Qa[0QNd[f;;S)CCP2M]F6ZRA_6RJId]UT86N5<Y(8eD6H/D;P2.N
// Y7+[)M^dXSDUY\<.Z\:,W9GV^c8@@TK\0?CEOKI^ULPCcP>A;D^J]KE7A:^-<J7H
// ,:8GgKEJ2^;IFa?-0(RJO(YJ9V9REg5C+R;#QT9=BU\-C_<,AW=/TQ6;4RHN_cD3
// ;#g->>?[b#HN,R>+KSE\BK/\<bN(##EZ\Wdd[,Z.cQ6IY-.(#PLL4RbSFa<7.19J
// 43PVF,cDbG2Q:0S=d4]DKOd?_@g7egU4=af\)7gfAZP]]J8U]K#N\Z:I-&=bVIU5
// _M3-?68f]N@(DD8Ke@K06bgT:T.,?OX#YaQ0_-K8=S+d^d@45Kcfad_bVEeS@#eV
// +SY/ObW#[IR?-\PgZYLP66=(15S2NSE_Z7VB204YY[OaM(CF<6<F<f5[AF/V<;0\
// I&2M.?a6D^V8YP8_-]0_E?77)0c+E9I26#@QN=?d)5]1\?,bA/L]^O@Y/(EV0:-U
// 7WO-#;XR:K1\G>eX<Bd)=_R&\G1NCgg2g0eB;#(]2(UK?XVTMe>D.20I&NV4;BI\
// ;V_7OPaN?#>KARG(1XX&^YZZE=EMD<ZU?XcP7DL3.L-U;(gbFXY_@P<1F58ZdBUM
// /7S__/\Lg,NY3:Qe;PaP^DT8>fH5@_6JUHc2NCS:2Da3MNODJ1J?Y-RVAeL6g?\3
// A8_+YA.5^P-S1d6=+1SS]c#)^AV/[ReD6@]0DfZ@Y#/1c0c_Fc=cI)F3ZH46]gJf
// ?_T=,8)<+X:9fX);FZ14(/-=+#\0RdFL,7b1SeeE1;GO\E6\V).0&T].bUJ.BDTQ
// ABE-TX-WaKJ&^b>?7^B429&8RWP+<S[J7F@a0dRSCZcYLZ&J,(GYQR)K,:V2BK>6
// D81Y^J>(CE&56QdPLVEecMFE;2)=;;6;_33BNR5]._-M.aWO5O)aY/(LW8H+HBLT
// _24CDZDF5T^31\_<Dd5/8gKF[2O<61WE4C,+3&OOMWV^77\27e@M@MK<RFIA5MM#
// 8BT&^Q\g.dM6A\UE6Qd<JLO:Y-S@8&a:+3ILb7;G>-Y:#6/<T4&GH^8;+C&9#&.&
// UU1c#gUMWE;._82\@#O+MYe9I:BIfe?G/I^>S<4<4gKHCEL0PT&WIQXQJ&S2e.-D
// QYB\V&IM5Yd/MI5E8OANDO,N\AT\K^PE5ZET[.NA^:33c\+AY>QP:1CFeWIP7?=>
// \g]C10J,XM\\818U@ZW?C9.5R1&g(<5EQASE)d9[Rg#TH13]K[[@I-gFZ7_&3_Ia
// V:ME=\JLFEK>?;&188E.dMgE)6]H8[P8DKNHN2dcN.],_)^c]d.(HMMb^PC_TN:7
// 73LH1]6.:b4ZJJ.,E?KB[3eV;;D=-4@.aPc8_e-)8D<(e(KJ&6O#Xf]M8GL5###=
// 1^XFJfAYYMC#I)56-#Ee]X,_4WGUT\>b9e6;O:a[gcdH[_Ye^S>CP>.Pe-D?HIUR
// \geLRX+C;3RQ_Tb&)=+HUWZA2+?R//VH#N82]#:df@]YV()_Y8CDU[_2;e)(?,22
// IDRP<Y318G8+Eb0_2:&)WWZ/&Qf/0cTIP<(8V66Y16XN>A5N?7Ia>WMCgfc5U^7)
// @6HLECefe3cg=Q8AHM\<FOITZ\9[(ADW2]VN95g&NXcY)Ng9G4fT2=MHZP84=-fR
// 5YPWM4(,R6X-CgMAN@VNJO-FZQ0<A^,U6/]W3DdXBN=<GgH^3:dN&J1(4d?(9PHM
// [b<5]FNL0?:)\fe>J(6Na+0(JU>CICPOZ.=,0]G#>eSZ.1W9K&;bg\U6-,]R3>)(
// QD+4PfMC;/]\JOEFC/626V1@ODV?2[Q_D+4TIbI4AI+,TLd1e>Z=T[edA5FN,OL_
// c:Ec;(AM:-831fc2c]X<90aSZ;.\R<P_\N;2LC:L/]]6HGA7@_5bU_C2)WGLI@\F
// +1X6UBH+?.E7/3_=.G80#R\HX];D_M8J)\^Y[?4Fd4+(MAO,G@K1B9IUYE>)^5R,
// =7]O3,&=A+8R^?41K_2OL[:c@Og^CH_<I_^HM:#cA++->KEf5@N\\C=)6N:g<+7[
// =A)#5(PQ,LS?3V&N_R]#QIJ#H1LAM-OTaGZF1.0BQ\6Ag<B72)MPDD&9)(I1\[Q(
// /d<95;L+W;?6K3\2:.F>+bXVVaY.C#94,\DegFF=NR=RMO-R(43<IC[JW8K7Vb>X
// #EgTK^e4UNRZc^YXI.\HWQ0+-+a=Q?XQ?aTJN[MFQM[I\Fd&4(J:f2G/\YP;P&0g
// #M+C:5N;NXKHe1cN-LH<0gI8,J+O/.bHXa,5+B0gdf3DCdAe/cBc^7P4H7CKZA=A
// @(W6cZ:2YKY[5=.Xd3@BCa8;EEF@dFY<CD&aF-CFG>#5B4@7d;3<g@DS2_QN<2)b
// 8fIG)G1CBNV=16f7(eE]&DNU)Z=d>ZFBX(>=Kc;[Eb6df(WJXMRG2[U4gLW[@MS>
// 7]g)HMdFb5XfdcC6ee>^H98G(+#]>H0DMJN-+[\gUE&P6_[F(#BH\[Afa&aK@Q?I
// f;(\/A+V:5N);.Q8(G46W-L&XPUGDEGB?N]@YTZB4fBEZT4B>\BR2@aFMFU\>P,V
// OC2gT6,a-+EB&P#W/T0Q98+&U=]R)f&R2-00Wb\g6g<CXcA-_eYJd<CITcVW>(WU
// ZK,DMBFIA/.d_81P-e=#Q-V,?)D1T+RBS/RRg?/W(+C:NSQ>),gPY)T73(KB7HT2
// JZJ_4&<f;7bXB+bXK<ZW1:gPU(:FR.=ac&5Z,PPOB.0\2+b2Z2_F=#QT@GMPURF.
// YP^ZV>NP[G:C1QFOMQ-BD7,\#VKf^XM7QX9PBfc\G\=QV))2.cf?\(\.HX]D_;6^
// EOKA=1#@D)XWVfd<d>^_UWQN1V-C2+WKaJc,Jf8H9:1_PSVCeIR2,>R@C#Q6=IKV
// 5cK)1OS)>CCQ2,=:<MeJ=(gLJY64Z&+M1C@cU;JeFJ>fA#.eaE.<>>e,VXCTYFGZ
// YXaC@^9:]URA^@:CDLfH?RDV5Jf+AIS?ObQIA9be0GbVAe6XH7:?6Q4I78\Y]+3R
// TW4dU84=P6>L_8e^L+J#-Xb=YW,5W)=J@-F-.5g:P[_=0.3YFN2#c8QYa0B[g82G
// ]a:cA2a,L3EPA#c#We#ZMa10d3[ZD#bJFAV,&PFNgVV_.L5R/4\[:?b;^CFYb/@4
// g++PH=&BY?MT5aH6.QPP^[WYF>]DDM-,d=FK&/^QSgN.7#[4<YQ__A)\-5R#:SQH
// 95F]BeVL9[UGYg>IHEG_d[D7Z^JDDC-HI8^_#+)dLGdQLa:<)#BYIcd]J94MH=I8
// THID1(P=XeL\JJMW4FGOgY3U.YJV7_0f3UJSNEg3GG3M([B]@^6[BKRHA:T2A\6\
// d@K=X?35fQIE?OO9abG94+TLH#7[XIgXJZZ\J77,__7PC,UU,)+??#ZMQDAA9PE+
// .8R1O6B,gUTR,aSJ]D+)-QgDaB]-(bOW40:bN,V.XOYUQ5+cVZ&_;N1;OV>46R2@
// MOLNNN)/L,3.JA(Y<@Y95TeK#)dA,8LXH)+Zf.VJ3bH-6\@Y\[2ALA8O2UGK&6[R
// T+2NA1gUOKTbQNQ(XI;].G\=Y8LV.LLNLRa><Ub7b+>-?D]5_(dcK.T#_CE2\]Z/
// .HCZC=BBU5@6&ZdSE7P]1g:)?C.CL?5T7<)_]R9)Y<-&PZ/I9gcEL3;A-9\UJc]X
// ?_@K]bX_BXBX4C\(;LIa/eEAc+Q.2B+NdG)Rc.-Z-P,HbN,,fP>NTGI)-OBXa@Ae
// VBWIMLaDB>cMF.[_Ga3DV]Zd]e/1XDeJWY:SI;Tba>E@5X=1DV7eTME4gJW0f?UV
// Segf1?-0GC+gbH9@0G(ddWP8?XS&IRfG>W:A3,SJ-30?.QQdK<?,\b8T<1cb]be[
// Z90fK&JI1@&VV?JMAa7C4^O\C6G?6+N^VQM:4BLg?JX60ZLU:g,G8JIJ>K4==X^>
// =NBa[5)U[\dASD=)\RXGC,_N?^KUa.]+Z.Y5gUW\Zc\F9MaXJW8?GJ2M\bYL]H9+
// O5<,>NOP;]B-23.:/^I.gGbNbG4F#9YF&QIK-fCL/:X?,(PO0++];@65\4&GS&Z]
// :,@J)Rg5P<&eZ=P>],(Q<)XfcC<O2&(REDT?B4?B6.BS9IW)1+9(Y8]Y2_JB#>5L
// U1>@+6FAWfa<9&2]LLT32+B^@A5C?Afcbg<2P6]0Gf>[=IRTDS&/2bdQ&&)Nc-C,
// \2\L2#cPOCQ@5+NFBUgdRHbBUP]Z;;0P^<=U)2G73PF2F[W\aXZX_(^AWQ_fA0EJ
// [GA:HFSbb.RRVZ];/0.aM,gNNNF4fQ6@.5FM;BeE;VC(>&[E4?M/ZR.MZ2AAVW=f
// =.IF0UQ+R#70-ZM,,J/Db;-/b?>cRQM<+AOTUM_8b9@g1Ed<J9UfY+_H=_WZN^fB
// 4GQDP<N..29:?P?)5&KVUFbI[^.40\J2V=O]VM8-_00gUc02L\\^XILG0f#FN:6G
// #2IgD(c=UV0;=Zd2ZDBJ.ORXYUK/O4VAXXG;Z4)YgJUa,/M<7I_86-@NcP-f4WR_
// EHX-3+.&<\U))gLHb+UTfKM^;L9)70OWYa,/EFDgX0QLXWQ0Y?EH>URW\fHV1B&^
// \&N7XVJ++EM)faH6G+0<NYeYdV&BM#W:>KcfS8M5c3;.MUF\d]PD1#IQO3&6R4V/
// [#Pe7YCgY(6K1RX8eg^@HQ&0T0(6a.eC-NN(f?YC6S;YXCU;aVfI_MR7JJVH\]HI
// 8DLE9+YGB>COBL@fSP)OOI=;J-UM(YDBHPQaK)1N=,&AITD:dP_6.dXILa#)<H,7
// R^cUD5+LX<;,&Te#PN5:Df<.bRT]MRdG8e5P(HALFI.6d.Q>3e5_Ma@BUQa>2G/(
// 922cJ/8=AS6RCJ&S1M_c5.DA(3LA[d8V/bQffV5HI7ECTYDLe>Y9TYLU@;DL2M[C
// Q]U8/6NM1+18L6KcB:<dPYI7:P7[OEH@L,bK;#/)_bJ425T2((fI9cN.RKN26+N5
// W+QVS4V+N/H>@NRW,7KAW[-4CTNG]VU=9Wd?PK9F_cf6aJCNf;NURO2cO=A;4J9S
// 3-d1(1:Xa/d1:4?+#2K@f?RZV[PdA)HC8;U4+&,>P<+5Jf)?AD[N((N-&D2TL9=O
// =V[G-M0;+MHG,(DIQYHP#>8>35b16.WU3<)X)7UTLQJ(]g,Ma-9W.07>FI,2F[_B
// 7_SW-=[D:<W0dGCGe0ERHV/-?ZaG@])\f(9CeCMbbYYHKZ#O)J5C.->1)g45PcKV
// 5]9;]6X-=DfWXA-W892(:+84/<PgM9BCX8TLOf=eCac6>M8<S@c[/Wgc3@T6:V91
// Jg2:32@-Q_B+C_R^Deb#cSIB8A9R1)G^4UG0=#]LTNB9G]33]5ZGO:I-&g\+3._=
// =4E+^f1&a@Y&/Bf/)f6@25.&;D61,XI?1.GM@65H<V_,9LTD>)a:/:O47RJ]B262
// QXCa,3/+3O9@ZF7[b[?).gE]>-.2,=\1fC@f<_LQWc7IXS]^1>TZU6.?KKMGXDR&
// 4^_2ADg^B[_0EBY(-8U1)ML)_AVZeQT7OaD5H?X50E246b^QC^N=cXFOHd4_HGe#
// eZPa@;E2+[8R],1E;:)YOC7(E0-L3M[TNK8T@R#AF.)JXHZE,bNTDLPOeL1-ZDX+
// gM+&OBba;VB@TbTGU#>DYaA2>5NQ)Q>R.J&6?PaB8._D5?+9.(_=72NI7S,7S+QI
// _L9Z77S+bf3CScNRIHBU]\g5Q4VM6GM7bETM(gE/E:_P(<ZU=A3/DN-=]I3Y(\#-
// FW0F39@VXU=1PB73:R(#1Ic#JRg)32a[,c4+-]E7NTd<1[11,JA&]0e8c^d2f5[H
// #?+(I.13RZ5UL3^O_S3&9b8HBP?6K1^&__Id@B5QG;)0=V().4<85[U>74.?Kc-C
// #IeDDRfGS:<9:O-\PH&5;4DECCG,=M(dTAdMR2;Bb\&g]#8gQfT]_##)dEW0HWBZ
// Q\3G/,&J1e0F=_YLa=-PdL>>(5;)RO.(=)_,CO2;2[AYNXR1TN5J(9bgGdCagLSS
// ef:YH[Z<<>1[O[:Pag42WAf14KMcSO4V(RC&LH,8WU7OKa;OSXIRac[<c=Mc,e1D
// K@875.9EB>-#)E,Q1Hdf497fW,>Wf_Q3.,?8YD?9S]O8MO77M./)02ccPdI6,42A
// +FG[-UAc6S1X>O@LI9d=DZ_#=a#WZ3e<<X/#-<]^H0C4+B(c<<c].]IT?fa8@Ne.
// A+SN;=6a>=D_K.5W>NF]/7bVJFJ<9WHP1(ce76LR4C7e]<2-4-CBKf>79BGF,ZWZ
// 7dHEMc.0S/Z6_T#e0S2+e^14K)g++)UMA-a]B>5G2\M7FV2MPRP(ZL39MBR2V4BQ
// 4VA+:O+-=,D5)VceI)g7;;-N<&J@Z.O.)-QHZJY:aVYBCII>UX7@APYIR;=+)?<V
// YL4EY?Wa[bX)cGM.#UA:0EA22bfePHZF3K\bd#P5:U4]#b(F[;VQP)\UJ5d+fXF0
// #<,3\L:EfFW\_[@^:R1X/G?Q9,]-gLL/68-B5B+3T//H4^PX\R#MQ-I)e&V6-&&;
// 5T,&CWL^[+M3.7E4F&.YYZGY^]2GAe\)_R[KN2=Q1N^5BVU=O&N75fTCLR)(NN0O
// RMc@_4)KBRT7GbUN@W[L@d<7Z.Y&FZ>[A?K4=08=b=e454Fd?4gTU@W-OD2:92/@
// DgF(c?DVGXQ7c]#)WH(f2&cN)HT+K.FP)TV<N+J8-Y-KWKQ1PZZLc^?)U=>+&\.>
// HVBOZV^PP:?OK\=\+d.WcTLO<ae\<.acM:0Y(GHNVEZPWgeSe.Q&4S/MVAXIMUM8
// aCG8YbB#6g6(O5:1BW\G,=/Ng#HEO^[a5.TPDZfOX7M8O/U8TM)7)f935#.TY/E.
// aaU+6_@McERXQK-=>7E)OK@CL;=2/T-WD3C,)IL??6;S?QGe>I2YIfAJ^3HQB@Z\
// :LN_RIJNB1E3>Z+3.UDdF,PgH&[d:935+c)-A38ZGR2-)<?]?.P[)eQ1J1e+<0gE
// ?W]1APg<AZa62E[8ZD[?@E]]]c9#H.HX)e&NP:95>AV=71;-YOK5&_S92W@+N_9_
// (KK1+fWK[)&B3OV^</Qb?PGNCWTc+bOAg[+K6)D@)ZLJXTRXKbH]XF.U.H<SD:11
// PQVI5=@eAN08=(Ie-H0JAODOYB@E1)2:=<0LG3#XXGd>A37UHDGI5d-_9^-9aI#I
// 7Oc:QO+UQe\^UgZZ)2#E_=B@6-,3E-:)8eGUbHA7g@SW.6RH=#R^If:Y6c[/cRM0
// ABHO=5U-d?+5Y,ETf89;=?\;9[=P#B3B=Lf565)gC:KGTT/>IX[D^_<>[C_L5E(3
// P]e[8^98C4^W1S(\S:V74BB@><B[d,W:/PgfJ&,bfD<//AM6E<]Na?V014WbJ-:N
// &b0H@6I>b_#KSUT4=)Z<#AXA+5_9aeR@HgBULTPQWCO6US.BCGFPM@L1FaTS?OB3
// G>)FC+)g,2=,SE8+>S-]C_U(0+f.BgB/#S>2&KgQ.FPF(W-.Hg]]0&@T_gfH>QMV
// I0=MDU/)::OZ/U&&PIdKdB1(@[A&Y243^^cP:,[PQPeI3fF@1KE&gTB&ZZ45<]_-
// <KU.Hf=,JPI]+gbc&2]e4BGeBNT1g@g8=?NC5]Ec]U0940D-C:_JW2&#CJM/JLN#
// =\B=b^9#<FYXR<J1gBKQ3Z2RFT&S@e#S0WFO,e\>]4fb@^T]E6agNYdVD8..85D&
// /E,9Zg0e\G#d>Q&dQaGf:?J1]I2\fe4>bZ:P.,02;7<M14C=^D7a8V_,Da5_R<b-
// U;I;75bW^UQgE]7SB8Bc=8EMSb28R9;g7,a6.C.B-:ADZ1TO=NaK91L&B>.V9Df0
// \Wg:,KNf]8_0&c1IBDN501-bcUCBWX=Ug=8T6FJ5;@7>PP+=?D&g)U5V3Q#/[Z</
// MB4<7:AKWe<eMO5U^AHFU>QR=AMa)QJ/-UM;/9f;T)C^J:E<RK9bcd-O>G5B9Q5f
// PK0Z)5QV\g<STJ];ZM2PO_1[803#U6Jf;Kg)L4fN2R_)GP9WaL5MF1Q&(CB4V5#f
// ZZ(;[>Q))?gO)a&\FH-#AeCW2:b(e-aV8EH_[&MX,BZH?1[(?TT)@9VRI^F7:Z)d
// M=()6OUF,WP/.D:.^:WEA3cXC866AEO?Y@=T=<DOZT8;X0[c_[,@KW\X4H=UR+>)
// F_0&M]8(D&VARcX?9>Y2H3egDC&.A,dFSA[+=N69+@>.,+bPXASCaP1?&Gf4b?PC
// 7XI7<XDeTW0>=2g@TK]B/#gP,dF/)YKHJ1Cb8CVHd(@-6-2S(QVAP(.-9\^W8Q1a
// X5#,1FD2@3Ld.bMdHYTMgX^bX]@IdQ8C60)X02EZULT2W3^#F:2IR(<IX^f7T-@K
// 8WL;ZMb9JUOD9<>\MY<0M-BX]4XW+).Kb&=]=G0Fd3FYS0a?7<4VA7(9(+<)N4)&
// a6XM]T?<J>P&9fY#Md:Z(gMbCR;AI7+NZ/JRUQfI)d5R&GL.YbFO-01Z<[H1a(O.
// K@cJgHI?1?C7>?(]=XX4.DRKaH5+U=D[3BR+K=+S&g><YAb))c8dG[X^WUI5ILOb
// 0dWX7aY]OO0YMdcCEGK3P27N]VfA0Mf3[XAPN+68XN=Z&=0Z0&OHTFT?[KHB10@?
// g3XP=AR+Z,64LYJ4ZDN0QQ1AKYYY+Yc^<.#()F_^Z\9U=HAK50^7<7S\[&S+(,_7
// Z,9PG\U;(9MF#SZI5+R\/U?<\C6[4fGH:#ZJFG&gAW.Z>gM8eAOZ4.1+Q]+VI>E2
// LgU[aO@cS&]K]Ya#E=1FFd7M?=3H_DGSMJ+ccBW<LU[.G-T];:>O8>B/^cA:XFC(
// ,O2gC.G>^-FaM[E)PdaSb>,<&9M9AXVSS9/eZ26E]VRZbb<6US[^PHb:M/Kg;+:5
// ZHYESSQO7a7N\=7J=T<aMd#\MXY0R/>^8,/=Z\,+M\71B_[0/C)#T)25EE/VaK[<
// ?B9-T4F[GN^g=e)?3LPH.I_F9Va#@GQ6PE;?1F)23AWd08R=P/dK2QTMbfeF/dX=
// [5LHQPV,X4H4Z^?_W3)?KV/)^<^5d(5_/d53?&=BLKgcPNPN&KcMe)1.@V3=NaTd
// 9Z_+=d_=J2K^^H2T,1eF5b;7&H,,LKe&HL;ed871OHE3b.C;/^>6K#]eAZS)4/U;
// +6FF1QCd/Oa4>:cc1Bc(-IDZ2QB(NVEDVfRAK;g\/?PS9EWc?@UEU(QF4TN(\Kb2
// fMI#T^043B/92[F012JV(\\&_9g\eD9_g@K-WW#]M2]3G^NWEYYDL<<I;O&b5@0T
// LUGK34F^B9=86X:16&KSUOLMHGL-4H.BRaM_+59b3VP833_\L]0_.<5#_D7)\LV,
// gS.YYV]?PJL<ONJ)O;)1_E0WAG@PZ10)&6Y#VeXcC+,4#B/S?0Z--c(3?1O5ZHdN
// :>EN,D5<ZYO?-SV#SOMcQ2M7[#A22V[1RCCAONM84(EWe_;C<aCC\YKAc/#QL&Ba
// K?M;FZ\B/+W.R0FF@:.,7)M@3D;9A:5)O,14Q^3N0WRbY^@2a]g\KS6?@c&)TEg_
// 4.[cCI_=AZS^^O-;G4Y/OA?gS02C(:Rd:ZH_UI/If-O7Z7Y?LHc^J_,L9_G.DUI/
// E3J&N=LVN_)3KMb>?+/-JbEA@bQ/./AabbH3X;Pc3,a.EeI,O:&WO0@L4US&^X\?
// D67AIG=?cXPC;-aB.,_-W^9=\.XR;#M6G.SeJC##KE^9Oc6g>OAOF5&6RFR#N()E
// ;A)I]FM=?OU\<AABPWO;=8F7BVbI<;g@+^JDYW45I3Q?K)J&4L1.T0HH.3ObHfZY
// M1f+X7N^^a.#(=,U1959gO/DgJ@bN7L3NPG2&J6^HSKH-#J)IB=K)8g01Jb46g2d
// 7AYBW/-+[GeP(#@M_?GYaD/g<^Yb>e50]EKcfUT#,=NQ9fb^CL_[17e70/WY>/c3
// ??-3S#)-EI?g-\Q)e8<+H8A[A]2TU.[7]X;90-1BCdU?_bN^>&P/6+S1bF]KQFE#
// I<fW@Jb;2bLT_PPbb>UFe042=5ggZ(=B:D>(_eFBL5]c6T/aa^D3B[Y5>a#3,WeS
// 3QWZA48Y+:VfX9AC(\T6a=,2UZTa3_D>OCG>;@4KO#=P5HHaF9FaeT-c6GH-Y;GZ
// :eOaF4<I)?9VK<N/eQ=-NJ[<RF7&&B6:/]7Y5@D@9)3H-P-Q=;KF.45REfWMdAOZ
// )Y&(]#P5(N:N):OJMY8&bSJGf98;bBQ<,XAU:eTY.2X,?]b[ZaLZHWSY;6P&8g_(
// >Qf#.MO,V2HC35TH?O]9KAa2B?Of]_>bQU490((<4ZUggW^BYg\[AB/YDX9>OF#N
// -,Z:I>)M2QV2:\R(BQ#MV<;1.RVRVa5eee)@NSEA087C22:)aaB?IK)8)H7RE;^)
// WM691VZ84-g_COUbb0:F#gQ#ZBES0L5(_2a0E^(&FO\OYSH02IW^?8Hd^I.TX]g8
// ),,+&D@._4/E/187(\C^\+2G\/D8I?4)BP<PWK#3BOe1X+.23H&:Z+LVaAgD3Q.O
// 9DW7VF3Me4_PZeW:+S[5X9D+-0X8&4\]g_6Bf;<J5=f5IB3J/^IS2Z+A<7.V[BNS
// ^GCIX16V\2S1Z]E5&)/WVNR]<EBZRW\]X6f9:=6<d,[<O/NFOIa\Y],+]WFYc#=4
// D<R/[>cPX[CKfL4Q_86U_&6XWJc)(4I_e7g4g\3ef7SO_RfY+F8TMFE@6HNfF8;(
// C)H[@?[?:_e@;1#.S7bgdEVbU.3ON1/)Rdb)Q9<^N:/[cC?:CU=Z^JYaDD+GW.26
// ME[K)BNQZCW^T9\64fYA8C.EGf,fZ]IN#RP^@BbD[,:BfA@+LHM@D,><Y_>dW+C6
// P)[K?W?Xb3(9E#7U#AJXPS6@8=aDE.?gHdgM[LM@7UPUgN#c.<08^0G&?Df-SBT=
// J03L71gfT10FeY+#](LM_+@N#gF_/8V&THXC+,5YJX^IJ(+<2(,Z78<IVBVKS\G6
// Mb(.&-YCZX>](\J_@NTH.,R4aZK-B+=ENY5G5T,f&Z5Qb/U7a5OR3)U;<CMUPXS,
// (1)9=4>_GV_\C73-55Oe5,Q,H)=/G0_TGI1=TOXFNZMGB(7N0aROOEFAN9J[.=/,
// ;>4Vd?^=U_RQf&V\61R:83^0\#0(P<4^J_edPAAfZ+=c7E1V5V4g9K3AFDPA,B30
// 1GYOJ9c,R8Ud74\E#<6U&2eC_EO>=H9BLb+9[NdCK9(@FUdL]9ADB]C.F#Zb2aA?
// :eR?:>:BM1J+]6@3E7T@51XX1CNTd\[]#L4e\B19gK9+AO:fbP7/W@5\?^=LB5K#
// ?>I^6_a#Ic/X/McBJU@WUc5LABVWCPg&K2&5cW(<PHcPQ1WW_JY&ML0&071@D6Ib
// a72BP[Ig#BN4b/0?U@XFYeBDXZ@=b:SR<=L7(ab(gGU.F3HX(QCUcc@GSZdNeQ](
// agO0U_5Tc0R=\?d-W3?W.EP^8]Xd^6EN^bLE?JI[c@QI]Z_6D6eN\4d#e6/I9,?S
// ]Jd:)2J;Q@<bV9F>_f1Ze8_KKFFJYIJ:DX@3E[QRggfe2Z0FRR)YW/-JF85Xf)V)
// T#92))fRa,gX,@,@R\V4Z=/2eY+7-a,G:I/]][KB6g(-9#YUTg3K/3a;eE)d1=I9
// Z55dWFQg_B;F<5BS1(G3G)2fDYN\TSaaC53JZ[#01eS;[9Ydd&8I[,<d8W+W)Hg<
// 179ea:Uf[b7?S2/X1[IaF.]g=]CLfO0;0XOf=?Ye=K3TEgHEFL;\;::UfQ0HIC+=
// 4@4CE+6DMU?R=V#.Zd0dQ/_[QYAN+VETYF&PW+P7WgS-#bLA85<@SII8^&[TXIOX
// D@8DOY;SYX@d7Y=D?2<TXB4ZB#;@Q2H1(8S<:c9B+;DGY1^Va4WM,/3#[ZT#gc5b
// (APba7HPe]LTKI6+CBP=;_XSEP)Q\NHA1@[=&E45=g=H;.4S]]aLN=?C<J^S0^AR
// 5Y]_?@X&Ib+(6<PQF7?@CAZ,@()[d\\84_Z4P>U20:V5HW5P8IU&>?S&,&\L9WVQ
// UKPXa7N/=Oe1QJ;O.C(^LAU/\_J?R8J.]e@7SI8E0L[-O=aW:B_b@NK.AOS,=?UJ
// g>;/9GgUO.B?CB]346:ADJNS(5;YS_><MIOA^_36UD0Q]@PP_/)Db^W-aD?,PP4#
// ,WeNZGX__R@<Qb::f&,45bE?K][S18=#Q-RRBO#QW@0H68b3>\8Z=J/b,/U.edO8
// C:93=00-3QfZVEGTI)YCF##Yb1?)-=Y/d<SIXgaUR>I.DX9_4YTaI042-CJ#?0Q?
// P5VH4cJQ:YC#_IRQ6E/4T.<WfO:OAELHAf,MS6e>_P(bPCg^87&A2&AK/W;#dD>A
// d:d&<S9d(LbXgEHZ[7XR#c)8BE=L.=)4NYRPW.3&g73?@gX&HbgF]cc&R,I2B2(^
// U^8F1<_(<=A6^;)XM<Y7[KYbKOB0?V<eX&RBDCP3:+91=#,-d(0GC:V-Z?UI(0fK
// >23/(bBa.7DGE02Z](a:\[6]G,9:0UGWD>FR^+W\e8S^#YFC1FM(-Y]&\I6Qe/.6
// =79O1bJeC9=.bM>@U&\g=,a\6/WSF=;@(e/bJQaEc7IXd_:#cPD_P=\6#Z_7;,(0
// UQ)LF&U>N+F_@UWd9S5?QS-JaD;_(0f;_@OK-YX^:S347&2BdQcW/)dOSc#f>6<B
// [>:_6X0UWYK2Q><954V>MSJ23McGRe8@NQC>CRH\5:+dR[TNEaIT6aL;d^a+@5N^
// ]?+&gI?3Z<)aTY_<a47X&.EJCA1UZ2d<@+FcWEfH\_DX6fAPPUTSAQ_+Td==.geC
// WFI^]7Ec@gM-]E5M7<WS&N?VCb7/PN(;BIEVY@2ZA5=R^7]&04a^BEP<@Fcf^TF#
// .V9BA[NS#>3#9VHQceOCc>?LRfNPVRQU<gaG9X;O(f<\?VA&8,V\@WO@Wd3<HEEI
// <_PIc)?A@eO];dfTJ[4XZ>TOA=19O5aaI;6<U(64;A5KX0[##OgN>A7;>IR::1.c
// 5T(_IP<VgU1,PeRIDKN^N=Y?:-)\8HGT69T8/aXR<\=c3]I(:-1#IE21>=FdW0-Y
// Y537&JT1g;aa&3U[\d.H)_ADg5adLbEDUM^PFV??RGAMY:=O]7[XU8)G?C0<AcU#
// 0],Re__3^4@@^Z>SDB&4eJ9eEKYd^SWYZVJb6b;L4R)&?^\RJ/cCHUC@O2KB/?>9
// [gV@Ua7P/GBJddFS<SY]XBHWK3dFR>1X^HJ2.AA9bU@_cT\&&,M.B#D/fQI=X8b,
// V,CESJ#ge^A3g8,;eGPCSZNgH,ES.O_HO)]>AY\I:Q)^5DK(g@#PY/;=G6+<cP..
// ^4DO?::\>@eB5c8cf>bJENdbH3NS:)7GZ6cCQ_N3OaJ(\,-EgC39FS9f_XN.\KV&
// dQM@I^ANT>Z:_Q7VG#ZH?3_=deL&Y&CdHAKAb96eGZW>I>L=C2QX)UWUWBNIdPYT
// KS6KH8T\@BUZV@eW43=]O>f\dM5IUIfV\+/e0TL)Ke+B8H?;Q?@Q>&D\]Q=R0b[b
// N(C;Ze-I0c:VNYC?JIY/_<W(>,Df[1#>(EVV+ee3.[==QBQTKJU0U0U-@,C-IW>Y
// /NTEg963.]F9X#5;))&RNW34,AYEXT2(S,H@V?g2+)^@JF2CDOM/]=b.+4GV@NJ=
// cL_P.b@aVP?^?#Ub_/M])-_>[#@\IPD^ONPC6e-<=BR/cSM?4UfAdR_1S;_ZPa)P
// \Y2FGDdP.QEP<_K+YC7[04?#+D9O,Fb;36N-I)0T.@[CD/bPgf1ZNQ4C_B@W)BSU
// 7KFZC/6.(/^dN@T>8E+.D@1C&Q:A\/1L-R]I^FXd?;W#K&.B&_5e47f#0.&AEe0P
// ,I/8=;#Ge3?CW.gW<E)^0Ve=GU<7<dM3QJ-^?V(<K#f3a/NA9c&J)f7L]GSFT.<Z
// H:@-^&=1=LW00^_SPE3d/4BFYO0RH+(7:OA:4H&O-\1SVd]5^9127>E5IfA.;AHJ
// TT7f1<>2)T9XYe&)>:_W>V+3YG9P0[[Q9NYf)-F:ce+ScZ32<?@E46bbAHU2O3LD
// H^)XHS1W#3F&4C:W^1[JWM4>VWEM]BRTEFWKe7(OS]RSc\OE[\[BaN5UITN=I&1C
// -b[QCVW7e@-IZCSHW4\;M(>);XWc]83VDCa#HgQPW5.9(Md]K3UQMea85H[-<<-_
// :O5FPf/]\@79Y;\[V[L(:b\39^0)#KG\aS49+)KY</FF_geJKMd_;).AHLH:WTT9
// \#AQW3B#FIe_.R(1)Z,@)ADUE<TZU(V,_c@;<f.^A]I8N1FB/S#HJ59aR4R@>KeY
// g8>)_c=5C_#WXO]=:ADPZf0f:eB1<I8V9BYUT-G]:]b1D=3/TQ\JI+[\:P&,Td+W
// H(R81>ADNXJ7:bI.7(Q#1>M=P+BA7FSU>WC87QMY/[P&#b]DPcW?RDHW<<0=LfRP
// a8XfFR=@O[W72NY0]3@3Zc>O)J3Mf\@X8\#^&S?\[MecF,R\T\J;B4a8#^_QUAI;
// ALb+\M98Xf6-NQ2<RM>a-FV<G>-NHW9=FQD@-=2Wf_)6d#E8,#66HP@53H+2841A
// JcLSaS?)[V7GOVQb^\3:cM^]H04[>_TI[Lg9>MXM8]<.MAXX7b-)_&O+H5-^7<?K
// T8J3YKSE)@+Tf#&BOfQ[IL[IPSdcC@Y=&A[5-;);20R2.54^#OC)8L/8V=g2C<T(
// M0_OYY0:BU@YJGERYS5F4GBCLSY>N5<)/;VALac)04dYIeDC0S9VW\8e#>ZKG[^+
// =KPZ&[AAf[ePJ^MOFJ]QJH^aL/Le9BdUAPe/.7R5BgY##;W1(fPJ/9,_+c+,\Y3+
// \-2(JKUP1a\FG)/Re9RW2SFP/BVWI=NS?C^DZ(FQf5&-c0F&gP(QSHBF00/]+?/D
// #;YSdMP+PFB==WB238)\^[cF6_FB_WdKOe1eL0R&D-^W<2BO^@bM4#8A]dC-V^g#
// E<&DXN9UWW)\VZI@0MX#=?<_DV<g\;^>^,+X2V&8;GM:Jge@6SSI8LSSa:]\\OQ&
// \:KN/1b-1de,C<[8363L_L?-Aa+>7fL7HO/c,+<>ZOXQQc<]E.9KE_^MdNFX?I8f
// @IgDM=XK2gLN&g>MBP>8?KCO#W(8Z.1EV0RORTX.->,G[^_]EF/PGLU(DL6C==+Q
// BX+C;>@AZH=e2[@=A[]0[cIIfd#XT.XaaO@C2Ab=4_;7JZ=(BAeKCI<J&22+F]b8
// ^4BFeW6gRMLO)>TO]IN7MI]]HBKa_f2c/Id5.fOE,8H]5]PXE>FZF_6]SBdV(+,g
// 71#5\)3TI]:N=N=1K/UL/fP.WV:a2^.?RfJ)R+-g&CEe2>V#b1&4WDHd7(]3.aYT
// ]9K.eGP9L67fU.T834fEgQ0(/2X&fXO+:=IAgL>#c:]_d1D;YTLL[(3O+8.G\H>9
// ::=Dc(PQUbL;.g2a[fT:ZfH\@a9F8^.;=-_2]?@:B)]0Zg@=dGM-N7UDWGfWHZc\
// R=DDMR,5ePUJ.F8.QCMOVYQd29(_Xc<0TEcY5X3Y6Hd[].A]XWK3RE+D.D6bSXTE
// W&CDIVZ@Ng;:541_agg1@cbOQFe(-G.cLT<;3N0SS2gb7-6e0BY[J9B>+g)?RM8T
// UVL_bBO\43L40D9@9eS([1&.D13aR-\\DIW[RK5SeS6QfT7G&CF2\F0.d_dM0gZ5
// AP)&fYeN7FW6/G_(RKWEd)Bf,1S:,@-?S\^2ND6-<P^OPFTZ],)U/<8N5\=cFKQC
// QB#<LbR[<\:=A3(T3H]66S[P?F8b)1@AP<CP=fPI;;IIPMH<#Wa8K(+@+=:d2XMg
// g@N\0#VdRV6.#FXRR#4XGVIZS-F_D(/#05GTDG>GQfM34+SVF3QYb)8K?O5D?F8e
// Y&gPfe6E;H1,7P6?a-QXL^Kgf-H;ZIf#5bMeX32@QT>eF8+-#EbbS[Q^V[V?fZcZ
// (X9OEg<S1N0(@UP#^9+VO@LLZcZ?.MQT@82^-EZ&M/OHN+a[H<&e[(#D?KMBd,T9
// V#RAX#BO@-LX82B4O)D3(;Z([24cK3\(0V<(d/c84][(M[=BN5?BAd=Sd2<DR0=F
// OB:1dQ+<D7C]TWCGT&b@Ff.6LD:5SCS:1AW5LC]b,0J6@/c-1,\Kg?0WFaGT^X]4
// EMbR1V(9\VR(NS</XedY<gf6a#NUO]Kg5\543AUU_&.[:7IVQ@c/^.B3PEbX]F.3
// KeT,=V(=BL5:/gf)K]-R9N[_ONV(2>CWWR.:=G8PSVV-:>\;O7NFB@QSO(]WI55Y
// b@E156KJ=B(ZW89FF;P(A[:>FO0eH,<2I_4)4N,NWQZKG2UNBK:1TQAZ;96WKMgf
// N#UK+#4Hc@0b(9c[.0fX>/(6;4d,T^OHWO7@+d]FfKE,3LLXM1:PJOcXT&G.,bY;
// )F_7=4MF8QZS9bF_6J3ITK@>RXJOU\B.0;F#E)C<X#P:aDQU0AYM0@C0PMg5(+EQ
// &XH<[aLL:JB2fF&a^AQ4-AF&0<^M,?(&ec((g+5N?#GM1)/5+8-dQ3XAZPcZOY6=
// 7?Bcg,=IIWY6//PR\Z11/0T@(.9f3/07ULH7E1F2QUA@;IB?B+ZXMN0Y6ZgZRecF
// P<CYK^cSZ_S/5DTA]D0NDK38[[cg@<:;+e.^HUM=16LF8;YQ1XeeaZWcVNAX?C>^
// PCYgfL22EOV?QFbU4g>1\&E\/@dCg7M?;PfcK:^&JgI4S#)+U\8?><RM6bH/I<6Z
// =KXKWgV7d;<P0PMF&XR8K50JcY3GNf]E4>L^d.H[fA,5+<bF9e-G7D^+cE8-Y:T7
// fQ;b?3ZR=ILUQ7egORNO3#0115)ZbZD,6O+_#?.?46Ca;ZCQY(WdJ<f9YB29<>Yg
// d-e?WP?;OT3>?UF#[PgGERZPa0&BR;c+F3/TSKgUQf?)BcDA]U40(AZedf]SY[W(
// :GL_EQaL-?#8\?#^J+X4@WM.-f:&5L\\FA@#UE+8_&AWOY;4M.XQ84LFQcEBf7A9
// S#Z+=66.c.0SV=>/#eSA,4c2H<R:RICb?F<:K6O;/EO\[UM-]N@R]V-];V>ET]<,
// LaT2fQHX-gg,4c.a)QP4b8D)-gCL[2QU-Z9DQ9<FgTT2P8ZU_\@=Ag25B,W/bHa<
// <MX;=;@,X8:HU\ACWdb+#G^?>]NZ+HM4Va[;C@8IWUa-2\MP3OL./f,Q9F&;[<HF
// eP5YSYQH,OI)Ee(J3[=6\VA:\@]T(HM1-?IbUG5:^6>;BSf+B+;RdX_)IZ5b7S_T
// :CH\8H6g,+55BL],gO;=dZ5Z1UT@;9<aDaK3VO.6=NcMU2-MS.)F&=U(Feg\U#)8
// ..VG;1)KC(e3caZI]][AaJ#6;:&[W+0@^1JS=C2C3I1Wag9QGg3T3e#7UdTZDQ:+
// ;:MPTO-Dd13U@H7b.4C(LSIK2E47YW)>)C/K<SJY6;?eF6>LKUdCcLFHS:KO4F[@
// F,FH9JIIC.eG<N\(78,MOD0c\L9aZY]fcP69#>#S7cVXX^=Z-M]O#H1<(1a,]VNM
// 8)_e49V5?HV+F3Y++JVAEJJATCg?V.?VE[O<A]QY1.@_=CacAX8N#A,QEAFW,.1M
// #NgEa,?29SH3)/-XH;dC8>KP2WgV9(24[PefcBH@9)\=gO4WfM=A7/5K]<XS\#ZC
// =P;U8aOSX9D1&JR]5#@7Fa_9^2BVJ5CNS#M7@aH)Wf>+F(Wd?Z7aV>JS)9\#Re9U
// <W\AgWDVOU+::7RJY=2+d==fAZ/EU/3LfLX.NZB0gXP1O>,c4-L73/+L@9^6X;\7
// =\2BEG<8>85:3,2RPW2>?R?-BLRLG.5LZXP0\#-3gF(F=4]e4I,UYYIGIYT/.W7c
// KD<S7KK@e[@Df/O[&FT2C1Xe6A,)<XZ)3#OX[O+=.Fa?IY7IZQe:g,KHXL3>+YJ/
// dE0G\IB7&J6N?e<<dF##T0fLE6I5^KR=2-6A5\P00Z(4=A_b91(7DHPaF&W5I-?c
// LAVEB>L.>/0FHe?I1e/>^@\8X[ZFLKJ:F@4#EZ[;?8]]A,9(+GKGPTYE#XfVH5/L
// V,IIQBV@2f:Sa.AfH\.UTZQ(-T-..0GUKY1WO4ET=(X<Z??Y\I24f9&(E@E(3a/]
// U\6QdJ^BY?E2QCN,2J6X5AU9@3X4K@Z<3.S:O;MIPLTL_>AK6(=+6SQ+?4S]>(]N
// :&@(CDXA823[BKLCBaH.VA82DV?1gTC2FLXY)+G?GX:J8;EVMf()XOg[(GP0]U&V
// @,e0,+R7Kg+68eM<UA<+LcV9S4c[XdEfCFPE2\E06bO1?^X:#KTOY6+_N@a#3>?V
// TL^F?bFC3SC71NagK&N-E:(Dac1Rbc\UU6)+,aQ-96T>)g(1,>9HX,:3S6C]R45:
// -^1L9(1Ya6FN(ff6,Eg_=3T443]LEHJcYYPA;(MbZKfLAL[f1KeK@b.SU@:bF.=F
// TPL-L,U6=V7;<)Q7SN3F[]SA?PAR6f3A+H)-@;>AI\GbIX=e:B@/(;[2f@3T9-\R
// \e=EgNLNG#[.MH26U7=]9EV>:4HPfJY-][U;1VG,eT,f\HG6&&-SD@AfFL\]Iea:
// HPZGH]LMfO)LL8Le@7H9GdDTF0TKP,.)_ZA6)8H#F>T)^0)Qg#/N]He&4]+G@23\
// 2O/9[U#;6=J8NbW9Z)g0=I]8_,GA]\aaAH3172YL(dF3R@EbRM>:20#&5-@]\-WG
// fYf]^baeZZT+VN.a[^AZV1N4^&D5QCdRJd96QJ?1X89,)df@b_f]YU2Qd,U\JBL7
// \;.06OL&7gOPG(M0I+V)4VA:0XGg-[fHE.TeJLRO#PeRDaOWDa_S[Zd4N&.)>8D1
// FS0?1NA)<:dG4fY\VK9L@#Rf4A<d)N(^IKF_YW)6BEK]RA[XDM^1@X@Q0CG:Ee@H
// eUaTL[WgNMCNVJLC+BB^UeLE479=6UK;Q)@VHNe;4A=aDC,R+#bfP3#OfK>JgH\U
// &>TV-HfT3[6/cS9Z2a7ZSX9W:]+WUaMB32(6A><G7SIE/CE\AP1#U0\G8YVG6DKO
// <H\U9NI]Dc#+]N1.;6&VW.)>bGXYS4^eI]9VW&cQN7TS^MMNO6dI],Tb33c\:MJ8
// F&WdH3&+C+O.E)>3P)^/8+PHd);+6-MIK9]PWf-(H8Te-ODWa^aCd>e7LgNaKDJO
// OUR6-BPH4=F02PJ:@6:MY3HGL-<?YBf]\E:Ta(1/A.&3+^fCN]d2(=Q5?7LZ@IF)
// GI0S61).e>P)9CHE;3FTP1W5JLO34Z>RfALUe3aKX7.)(eB@&8BGM;\DW1([=N_B
// ,-_Tg,\=P:EK3J=.X9PF]7@UQ9e]X:H&_+LXNA8.N>K^f](_[#[df;c](O6UE_;F
// Eg+B=LX\WW?#Zdd+-<ZEC#PPVKJDH>+Y:IM(,aR&/CRQbKLX#BWT;:fG22)F^edN
// 9[M\TG0&QZfF338.K(NBM-9LBTJ\)1AB8Ne:K8S&_C?//ZCd<?YFGTT2/.]6b[O]
// 9W]/\Y-1#HERPV#C,/b[Bd4f8O^^>V&[N8#6@3UZAM=G5ZJLI@9=PO7U,L-NM8[B
// cOT<>a6\<@U9>[XM_gY:Y?NCJ]NU7B0cKG?b[9:G\<BH4dR_e)14BD9Y6\IY-6NO
// ?M&0^c@8d^60]KcI=Od<U3X1DbTU4J;e9K.G;4\Rd&9-+RWe\4A_.>[00N(V1OEP
// bK_O?/S3P0X9.VSDf;&&2C6T_1KWfHK^8Nd^3+<De+bKEAKK,-FM1EPTP()fE3NI
// eMeP/:7.cO^Va>3e.HGa^K\b8)7FRJSSX5L-XU-b]T3;/0]Bgc//QHRJGGT26XWM
// 0@QVQ_c-;A<.\Q-/YM)Gggf,VO+d2E?JO]K;C7,<-]AbgO9_P\[,CgONZ0\K)Qdb
// ^VN9FW#aF)EXW/gC[H)?3N,;@8fg+BRbIOT_UM[LQL<241HNAg@HL\5McM#\=MW<
// ,9#+YPHd2UE5#C#_X?f]U=CeMc@b=@+(IN@,U5#-HUcI0N92HCdRfQWVF4<[1g6[
// b654UFOU-80N)M(ML\C1-5XI&1[bK@E_[EW14U(L.B28YH.KTU,E87MT8;P_QIgf
// ?JEA#-bSLV,V6P;K:8+@[(F&JCS-@^dMVA7OX^.P:g)]@C#A3R@CL^S+-^&TPZ-S
// gbZ5>(YeD>c#b0M.bf4C;R>1Cg1ZGH?,db4\52f<,]8M8))Fc,P9-@&:bL-6&1+#
// A>&-6a:P\D3e[J4[B]G8^L98RRaM(DbBW.#L6&FO93ag_@?LI7e>A4b.B1-N9;)V
// 32L=B<@CLM4W/XUK<>EVZXJH#R9afM6.M#G+_L75D#2aMBO?>^g?^_3M-U]N=c_0
// -QMgUJWQ/b?G1D]c:V7Bc51R)EBU0d-OUY_HC..4Z//6R^C_(9)facGcS-.3fY5F
// .),[#=Wf_6[2]SYFdaP,O7UagAX=PPZZ]U.>H,S]&2?Cbd?9R3M>(@QS48R.D627
// [LB@.GJeLRgFeTdd.API2D#\^#_6BJ+g00cW^M^AIbfN(Z;(CgT)PO0:DI]g066/
// R^2.9)d1dMQH.a8f0Re0W]U,RK\[LE6SCVP)/d,_Q>?0WTY1#fB\PRS)]:M<g0^[
// +b#&[,J^b[gb,):TA>W=(9E,HN]/N@_&791MJ;&>,S4:AN)GUB^7#Y]#)PfT63O0
// ??P90&+a)W3&13@3DF(]MQXYOGYQ)2df=+;HY\K]/.XPZKCO.U)8MU/Q)D:O.162
// ag74ME7,B>R<DEX:_#QSS,5G;^+PXM0RBOV<a(Ie<0WENQH9[f4=C1T.KM54@HX(
// ;?0e\HY1FA6;;dD:6ZPe]<bdcY];QMP^0IQ)^f6Ja^\JXOF#@/a6/Q]8Q@3,+ea;
// 9(8)@O131JEf;;K8bfc&I5?&[Db\IF+G\IWU7<1^Z&.3/:7F02T64A]F<1)84U+g
// C6<@#UD1?1)-3(1TCY1;7GEBcH+O;309\NgW<R<\I\:MfUfDRDR\@8G\.,[:K8E#
// R5f&_(HJFe3JC]>\.Z9E)=C7,SHO=+R06149LGGQ6JN3&Q8.UUFbGV0Y=YW/B0:8
// _eRc\P[\#A60FFE_/7TJ/75Z^F,76P=dP]6I3#0K7]KF9#CdVA:S0FG@0?V8(?-b
// ddL<=b+.664WT7XET)==8RQXPTRHB+DN[OZ9AcTX_/:_TgM&&]4G5RRE:\J678/P
// T.4H+^JH<Ae;C;<O6+<1O7SKLDc]LdM\<3ZC[#]KM2P._Q+Z8CUI6;_B_O5)E33O
// ?1E^CQ7@Ia>:b;W)U2.Pf]g3P)G;WIQ5?\eV2^W#PX<?\EgD->:_e02GP.U7)9(b
// >WDS;/;(1#VPO8bE95>9G>(:0AOK5BH@\8<8G1cU1/PET66[J+]@(XAe>TdR@4Sb
// ac#\e44d]bd[:D#/-I-cRF:^W39:.J=&)3NEX2YM3]F^#WG&].2d/;;e7>B=J(>V
// GKT><UG1dbfSc4e/.<:MZGMU:[):0>QIL08WCbL_/ZdFCIY5?K\f+a+EFK8\K-..
// H&BbMWd?Ug6e8T+_f@Ia#)-U<,,26W,0UM4U\Fg6F:DK781NaD8Y(3E54LRd8[MG
// #-]L)]5EgYNUYGS(?g#KJ.W&\0W:Vd6V?^HA=S,JL_W\Ag4O<+S:c>gZL4:HE1e#
// :^-cI+?16SV8aIEAc,aODT\\[LA>&TY25(F[^Fc#Me?c#^=67#GF9,EY585+=L)Y
// AN2KTLQ@dJ2\)f02ZcYAA7cI_^<X7C==811ffD?]XOPK_N_[aWBGH@C+H>@(UNPS
// [1Y5]f3>RFH;S?<A@D6#H&XNLEF.f\e)(:T#g)]L46#FDSgdcK#XPQ(\M.Ea+6BY
// ]PN_[,]fHS:F(##H&TdF[Fd0HaGOYQ=X\dTSe#/S=FY=6=>]#_fR5[,H1g<F1L,Y
// &/YO]WCQYUK2HZD)bg->4/D;DAY(/K<eM#=7>6,X&@fAO<C2;/SMO\SeW]ZXZYH[
// NcO0A<(HfBZ)?J>9&a7FTAPH^1ddTK#\GH91fW^;Y,-,Oa)>dOgJN[7R2CY=eWKT
// M[B8:I1M<UJ2);I;G:d/W\)\IId)([C@=f(TYJT_/E4FFG,LTJPUC^7/SJJXHMRV
// B-5DFK=6N>6D5C1QcT^KQbaPONVR[(FO6:c@E=c5.Mg3.JDR7KLfYC<Xf:5RU4P@
// (A\Hb>OS0V)85.UFPEZ7F9[XJcORTLV3:M]cRVG^F\A)eSA)KKN.aKSH<^M0#)2)
// /Z,cGWc;RWf^QJAHSRZPZ&We8IDXF;GfH/(8[cGY@,)Y]LWGLcXN7TEZ+f+UMAbH
// 2@#68]D/_8TL]c0OY=RI/3>bAN@Z,]<d]P1-\<,cU7CF[c.I5&cXJKgb_Q7N;^@<
// 6+BAeY_0,PObf4VX)\2ZU<ZLA97_14eB/Y^&JDNWHI)P&)cQ5F915DJGc5UAb1Jf
// e4;PeXG=WLSFbU[SL9_8gKZ5d0Rb,7)MDFI(.PbMSd1FTJ20BB)V#2bgI7SEWfe7
// ]<+c@;J]T6^)=&X+8(0aJ8.EHGVGFT11=W5f)Z.GAWW9S:/@W_G24d?3.2cD\7SI
// #SLb#:&V29I[&#^_.5I6bR-(:^S6[^2(&QCcJBCg:aUXB:G>BJ?KUN@/Ne6EUJ09
// WXaNSc\2W8;5X;R2XCNWYPcA3G_?J8>#Xf^F4.C0f6#5TPB@\(S3RD.Q9?ZVF]Da
// ggb1XX<I9fdT];X8<36_AA(4UJJL<^.+OeN@R_fK_0CH57XWd\HRG-9gcLa070g7
// ,4FJS(4c;N_&=c,2BSH2HefT?-\N<D=ZL27+07@-_F>>YCaA)_#Hd_HfKG3FKP,S
// Z0(6OK]T\^7R6LK17+Q<OETg@]IA<94I20]9LR=#8GC-N=@>U]V>#=_FCe\A([E-
// -KTOeMca8G6X4Y@8Y0]<;9M1VD#&eMdg7:)N2(0M9@5g1dR>F3[.[&g:V3Pc@Dd2
// <M2,Bc.#eE9Jd<LeB&f=[)R6J=W8/dE#>KD2[VA?4aagCBCM#dEJ.Z-J&0W2UcD/
// ]8V\C0TIcV)fE#H:bLI)X[QC8KM&OWg1-cQ4V&d8-L2K>e]][M)fTL[LT&\.SVO0
// VVBQX>V]4&E.-1OPNBG\^,NH<6P&#g;^P_WQ\W80,a:/QG?0BW7M.,CbJaD#?UN^
// /&Ee\9XJB5?JV#LV7JA&2MGJ,eW;S]62)?(MbDNGZ-(fM=E>3>[[=ZECWZ9XUU5?
// PB+AccD:9(S/JaT5aL1JcY35,45Se41bA_:D8DQ1W.:8\<WQ/3I1S??YPTPBY=^V
// 65f3OU=/G;^Ic0(fU9S7/c/AOWeDR^DNB,@QMB0S-FP5e\[3dM3LO#3:bdZR[2JE
// ,ZO@FRTXVB+P+(9O[DfT9ee,U-LLdVCS08f^3T2f_cR:6CN]>NCefa\R4G@5a8&F
// /S[d6fgAB2(EY:_,7][K:L3=>=(a(O2JZ)UF(TKR_E+aX)&N/\\46&R_]?FaPDUc
// eZ(O\7c^LP&\1e>&[W#F>4+_ECM:ZB#3>PC4<+e+Q-@BX#_dCF?IKU0f?2I=S=>V
// >17Wg--W\a4YT(&4=Ufc@+>LLXKW^/3EPSII.S\X/V2N-aDU.H]XY),=@\fT9(S9
// SQCQ_a\Tc)Z9NVdJAEZASIEg(NZ.NF90JY<LJT;XVI_VJbG8Oc-FOfQUAAS.Og,(
// =+WPb-T1=WWb1@Va6&&/3O=>L)e;WP@;4:VFN1R-d?FXWPPB<b&A_C6/EJ#Qd4D@
// DOd>eJ@TbX;e(PE,S;G6@:)7FOJZNTcPg2[^dTU7dO(D3[.T039,)_a3(MMJW_;Q
// _/9[,8K#ZYPFU==/7OD59@FLZc_)YY3TPFZ^J03-FD7T1,0KX;W#1W.L=>AZ>L9W
// YO0S;NF&]M+RH@73Z&5E3]aCY2UF)bFO^_(B>3e=RQ+_eX>9>K1=fFd>3aAR^LX-
// QU>I490C2DRCdc4b&YaTKD6K6-A,)E[,#?V1/&3EVc3c<(7a7N])T,]1AI4B4:_^
// (6P#MJgJNeXgX0^SR(8+N-7#@YI[=B1Q5/XKd5Hg,fLLe2E534T\3Y2FfSa#6L1)
// /\;?E2+L3)LQ_XSF;[V7T(^-VQK(MdbTTN^(6>K^XK<#Fe3=Z?W,V1]Z;UL-SXf6
// O,W>-?N_@NV8ZV/8>SNb4Q_I:161g?aRM93OY/G_g?830)cCYRBZ/S+I#F#UFTOA
// OFaM&1#ZII@g?.^0d/M[+;1C0479bIK[[F)I@&^U2_>YKAdSa/Ic8R&EA5>-&(fC
// a7F3E0aBaM:8P;=f_1\g;,.geQeZQ<aC4+f4WA^N2HD83KK<,8g[VTfAVbM7YKeV
// ?&,D(H6^IO?(+ON>]AD3]>3QQ>>0CX.#YG.Q>MX(,=:M70R/&#KS\P)E=B1_ENPS
// >1YA5U3I,7)a,J6+&H/,gL1</P/PGS^4I:8FC5_PXV>J6.4T)0K3//Lg9L\fVVe0
// &K(L]S\Nd7Tg<<V0EdcPHP^+KX</][?RgSHfa3GZ-(bH>>aP4abB.=&N>&cU7932
// ]KL50HZQV+e6eT^ae5eJMe5?b,B=QH(E1EN1g59YHEAT76a.A&R-X=R>A>PA9b9Z
// >C#c-[82GY-d47ae<)#Q3cALV=?#bV<C<I6#M>e?4Y8:VM/UJF5YcFMe,03F5)^>
// ZNKH1:HDP6:YUS[e<3B\Q9+H^abVIH_[Z_)3MJQ\[-U]V6SSEL;/R&S13WV:YT7-
// _UMeE,\KPb_1VT7:5/a^I8[eQgf5RHSWQcF6I,K0+[e/?,89UfGLDdDYZM)1#I<;
// 3T?S(CC)Cf87a+9@90:ENTUZ<R-aIUAeZ.W/[/@c2FX+X>9EHPK5VK7EeQCdc==E
// U#/6b9^P(XTXH(7)63Z3A;2P:1K#DMQ9QKCLa28JITWIe7R=>6EM2T>0[H2CU-AU
// ,Q>1E&O_&2d6LBfR[Y(.N+I/@X(U_#<eKOZKZVI0/7@8+U;SdJ^^[2EdT5L1X7K&
// VESZB.>>4=XYM_bLDBP-B-JQ:#?AQLaH=-RD.QURDMeFbdPCd4M]70e.SC;/#8]W
// eCX@8/&L>Pe^ORC4(M9dV.6.HQeeZ88;&=W<_J2+9-c.5Y>,#D1(?-)/#LV.W^RQ
// G?VMEaZ-GgL(:[XUbZ8K]0N3d4PY(MbICE1D3&<OT7RCE3^E?0g;..KGJ_bE^FVK
// /bATcfG-_N6aVZO6KQM&DBC\W<\0HZ6P85;N=/29DTZC9O&M:)D\B^dYXE?+A^@8
// 0KZ#/A6/a:;dbY#5]F(],V37K03bJIB_DgT;0^&XX:13[?Z7;V&f_dTIOUU7_3dY
// TIg><g@I?K++:9Z-HRW8<fYQ+QW=4BgK=>C59VX\O[D,4WefcTPc63QfI\d0Q<6L
// Y>_O/[)]XES&(PR\:HMUV\Nf:YPW9+76^J8,RA7(F9X#TR,EL,Db:^@MZ57DcC@.
// (f#^dRQfW<d1[ZE:/d?GTR_]#@6KZRG]N3:M?J1_S1NSSGCddE5Y37]CHSQ6YUa9
// 77AFWYM#W9(cZ#ZI;HU4MP\PVKA4U5NCKc9I2FH:WcR9;E]62D_eR?<^VTX-)d+Q
// JGIDK\AN90G30NSX,PDWRF5d1/f38\CC6^Qe_(3.]0F</G/S9,NEOAX5>N9\G=d&
// ]R#.ZJ#S3D#c]?+K]6eK2^eMW)\1&-]PN<\<M+O?E-V?U>,Qc6gWARE#7aLYCQf,
// M-\:6V0fD)IA4b4<Sg@Y#6/+)+WH32V_Z2f.6(HZT8:-1BJbA[Z9R_I;O?[>XD&4
// (eL[5=W^aeS5G&8I;Y=?Ya[+TC_19&73NOT+43H;>6G6XJ7&,KLG4_NN^fXOV)MP
// f)6Z.SBg;(c[@U=[6^J:J8>UbW=fK<I#3KN4&^Y:OXT,998QP#IGXB2]OT1ZZ=]4
// ;47e2Na&>d4CNJ_aH]d==_7(4KLgJM#ZO[;>O?e.HLNE3Gd(:EX1b+2=NS+eZH45
// 5\RVcf=8W;<+U@3?1MF3NgRFN]T;SQLSNY#UNS>V@4=Od1=+:1?]+2/#]MY=:PZU
// I)Pf9K,MeeC0FHT/IReQ#PZ40eETA7f.QQ14^)=R<ePUfYW(g2<MY8G)@.HR1.(R
// 3/+EH]aEDP<^I?1JE?;5b>egH-DFQ.TQ(>3+)L;L?-NS+MH06NQ?GJgLN\A\\6JI
// UM-PU2Wd5DM[?V.b&I9HE-/?C,=AdBX#dONSPBVAH;/VLNH&UX6(gCQQ#3@(R9aS
// b(IdL=V&>B=98KcF4=Q6a9cAb,V=1AZfXf9G4LS^^/:K3I4G:,:AANSa3FX)K+bV
// /9/&JP[]N4@E#>3(4Ma#E9b-&a&^>[f74@Z.Me0R(]OL[DMa<0ACR.bNG82J+B0T
// +?8V,86<OW61Ha:ZCO8G(JK-L1=Y1JECC<d#(A>1#eMK\^FHBbR:3]B,<]V6N].K
// ,C3C2_D-^H2_1W3-<C5-\O#D\:#4\TDbAB;3K9=a@Gfa-N&K]eB9;@&3SZO@M^H+
// &]BBY/9<O;HRAZWH?/^N5:3c23SA1?/gW+)@E<_f>+f8)N-16Qd];405/;\IM#8&
// ?c<b2<b4BQ1XGAO8^6T0MI6g48Y[9?_G\>B;W2[Tf=9)Rb=K&43US<4>C?;K/(/(
// W-]D5f0#<O,7RXK8050O\dgbI_;DP7B=fV8U[=.d9G3T-I.CO?.S&7&5+ONDe;-=
// H=M?M3]OCD]_C]fCE)UE@9.^[IF]].3QTPScfYT8Dc<VLD7RW/W:d?A406e46MZa
// S]fY^dSO8c;=&G_I-.K0R/VQ&[:G&W/)NK@gEU4#3.#JZ.J_d8QdB>Na&ZZ_bSBC
// BYaO]0]f8DRf\UO&Bb=I#O?4(MXf6E\,,9KT/5OV^&RGO1JL(XGM/;-)KWP[e)EU
// P54&Z(A>JYU:#_<gEJV/Z7LA\Mb#b#<4/L\9Ta_b?2L0Y9b26X[?V9(TOdULZX?G
// <JS/PSPWGS8Y@+4X,XJULRL.HS&SDVg=@VEaUc_Xe<dD^3#aP^@GCb)8I_4Td,2&
// I+<TQacJ]=]<(O)>6<</[Od_&7O]-Zg9KP@;MCcKeQ+E-32A^FSCDe&AIMSEZ7U_
// @dCA3ANSM)32eL?d[X_[eHV<)6\](JOC[+]GF9<gf&4:TKG9:IbV&EOa(@5SfFI^
// B9T0NE^]-Te6,.7E^2[Pc=2UC1W6E28:#2EXLb0ZNRYSA?N[+-cSea39.)9\W-46
// 5O4[BK&LL,VN>=b9(4^7,2e,LI-D-TQ)(KfX&6T.fB97J.aV\d]@&7U7V7.#)-5\
// [WI<G6W.8RU]B-(_)#T\cRGA6&DT-2Q9b<ZMBb^Dc^)4)/]N]8:SXb27;PDd5YD[
// -fT&A&G;<4edf_(;]_fS/A7:NUQ.gOF1;9@0@a\>7?2I#CD(gOD<WF)#-fDaJOJJ
// \1V4:+@b92&?2&T\\W@DG)P1P<(?\4=[1O);N1Y_^IVbfN.7S5N(-Q;UaM+<?#J/
// 2VU#>K-J][:PW/b.)QH3+C<5^:B)cMH7JH[\R_C&=;VRc(:F^ZVYFFY89_G/C);a
// @PW.@Y295D+V0?H5@1>Ec[DFC/3BNDDIHKO5[A&+CG071A&Zb<[ecXC]g50=8<QG
// GVJJ::^N_#g.5a:@K.?cT>Q2.c3U<F:DU&-I)DR:BH1[2G@<B)Bd?&CP2[F6=365
// @U>cC96^1d)(b8VU31XS39)=++JMXOYMJ-:P8ca6CaV9IR[AMEM0EI>RHY=O1X_6
// ++C(XQ(GOI^3<VFM(52;:^fCG89R.a.AZV<EVd8,(<K@AC,H0P?Z8gVR?E@RR-DU
// 9,>EW/1G_6V)X<2-Ha:K&gRZBVeOU),Mb-8AXWR:J]_Fd+/;#E<f-2W<JXE)be:2
// fgIf4NZP55L@S=(Ue+E^UgV&_8D]MYOD_#3-^R0b3T4)?b@6F&.H=84F:@+@:08F
// cK\KB/\X0S;<5IG;N.0+0<_c,+.<33cSA/&)a4L>BH),/:@d=;^NKCgVPe_;7H;e
// ,&Kc@1?]dXK.bP6>V<DLQY1B2Mga?E:,1WK3LEJ9aB(Q5LUaRg2B&BI#7-RSH2R#
// Q[W)f5DC7>)KQ@]9O29-ON]]92_eI_H)cE/;g@]-OeR2Q+<<#@5Kd0gX@?]Y@_\3
// P+Jc\c:.-Y4(b,]YA&,6-^gL1I>(.WS2JGR>=..6GK\Q,NL;f\MN7HNd2g:DegV3
// >3IG46J6Wd5YLd&J2RVe9b\5#e4AW:NeZR7+#=#B.N2:fVW[(aK=QDSK5@-(^.2R
// H5dQS9ZL_;91&F6PgD>NW>g0)K=VT?[QCT3^c\4X^fQ;WAa.A@ZWKMMWg3\9_DW@
// V7XF20YNg(/9OfgQ_-aKH9[-X6^.eJDVR+#OFB23LIR7@[cVa64])I?]<.POV9L:
// @fR+GRd(+SW3E?gBCI;g^ZB.?YK=HR3eEZ#Vg(8P_b361,=c3-R)1JV#(4gPX?R/
// N<MMRJLf_:TTI]KNIRAVU]-4bN>c_,.6,Fg8S8R8/H[-aS+N;<^DeC,3X2^KARV[
// B8gL3,1FQC@P&)BgO>Y5AXS_f=CgDUTG_Y3Hf9a3,=C/?,T2SVZ;NH#F^&L_HBP]
// HA)T6YZFP32eNF@+-4K6=AARH#]&9HCI+F]0BV1=5,?fNEW90F&N91E=4S\b=8XH
// C-=W^B.3+ORF=133]T[AF@EQ.M9T>3e(K\\MY-C/YQQ7>e0A,>+F=,?:E;).RW0I
// \-7#dC^GMBe1AUC76?DF3S?EI(eBY6fVS@88[QTMDc]c^e,FeNF8Z4W0Q@=3)7+V
// JX;fLAT@Y^_bDDCQPa8W_]@ZU)1_0MI5H^f)D50F4Zf,Da/;.ZW=ZLMCZd=PS++L
// 8JB#8(g8g81-NW/+gX5V(=,S9HYY#d\KAA&f</U76&cf(47De1M=1WNFP8Fdc&ZR
// <-#:C?7L@(?YL,SB7PJBH4E#THX<McDAf8BR]bV8e-8HW&MYBV-GUS8-fR^.VXB(
// K)FBW;R2+9/YOJ+#61OPB;9QW;U).\1V)HLWR2D8;Y:7X(L/Z=<:K#/c4LCQLTYa
// )-X1\VWIM\^5MM&9Q_6?W(=EF8Qg&d:YTI2D3aXJU6VEXKb86T63?gX]307A98@P
// dS2OB1aX\TX.Tb1Rg)(P@,ZU;KgNY^2e.&JMA@5CC[F_Bf/g4/#)NHBXE&0N35>c
// 9M7Ab40#Yd]L:VTIBR7]W@/TSaVHSG;N()(Rb0)(K42=#>+Q/>GND;BE+0Z)OXP9
// HBS+NIPeRd?KQJ&IK<DB^KHd@;/@Mb30GL,da^Te;_+._X:6@Ia#1>]AGQHUDbg(
// ^CY6Je#SA,0C9#KWVQgIYC?R\]Bda0MFL]_I&3C&LHF+WeV9.Ga6DW9C0.9g-//)
// QTHXA\9)=N3dZELZ<MHW:Y4>O:6_Sd(0CY2-1@2g(>C,Aab6BV.4#aPQ4bZceAR6
// d9(90Q\]:CBOF?U6MOQ\II,2?<)[1^@:<L&aN3-_56Le33EY9#-Ob0JY-^)^KNJ(
// O7]&@-TYC\/gAQe/37.WP1X\4+@cES1][BX\,UI^KD3W9f<Y3T00#GBg)Wb4ZcYV
// #8MIVJJ;(>O3Ead@QMS(HCfE<3a^eGW_9_g(,gT?T<bQ1/UHT/(e/SY+5gAN-4&?
// IL4bR##a[bLXD&eA_c)Hc>C20QSW?Xe,O8b0NUcYeE&b[gd[BfGPGA/2_KgMQ>A,
// 8e\BTNg3:1]F_]f\-PLX;ac^V&a[O;G718R[>bgLQ:+g1Y]WRe_)P280=.g]S/M5
// YT6S9(,/<a0=#[KIED1BN?7AV0f8C<P63LHOdS[(6AgO>cLQKTB]N^[6._.3L3V,
// M9USc2KH>KGNA;M+XN8)P7C;baV7fYb&b>4=4_75W>;X-JI^G@IYX]EU;UaC#_2M
// e,[C&W(N1@#BX,VU5+R]2<gHdXY.T/dWU>#9OXUZd?gE+?#ffg?M4@=UL0FXBIKF
// ;aK(=O#:JEUg8JN-SXP1MI)c5Y8Z?ESeD[WQ-S[Yb?R<SW/C=^[J0/)@<Y_T)&W7
// L#aPZW3Vc[H-DaXCDd0;fDML5#4ZBfXbO-RZXW<Kc6;Yd]5/.e#9\UBcRGY\W@C/
// CN79Nc>82,01[:E13H9W9;M_^C&b;c0A<_L?1S[[;)I;I05@2-O6<6PL:L@UA<&S
// W\];LGc-TTGDdMTbX4(\f07<cD)^M2T8#.QcVF4Q-a]K_+_TfebG9b6N^TQ5K]ZG
// K3(/CY5SSOF>LZ^d]\9F5)EFfW6N)]g)>g7MSF59X^^G<AB/:]?K?+H3YW6gZRS/
// 6S+)6d:IJLA1#?cZ:X/DHK439]OVJLXC]T[Z5aG>7..XQ1_Zdc[0L<>@\SHN4SGK
// 7YgSddP0=KC_Xb+c7JeJU+K@K-B+Xe)cBGTK4_3(+NRX/[NdVfbM4I?Y+b3T,,<<
// ^1Ye&b0cA4YF@]&TZ-(-0cR?YRIJ3/AUMHU=>W,W:]EGQDZNc3XS;dPK.T>Uf_8d
// #CYK8[daN3gCaSI<=B+P<W8Tf_,0dMDTRFK?+feJ7AHF;[=?.e/(:]8<fAL_bQ:A
// Qd<1ZA>/VgMBcWFd\5MO#E/I.fNVa3/K/@W#5[<N<<T>Hb\6a6P;/ULACV;/49(Z
// <025#+V#>0YGGAf_QA2FQ;_f2,(O,-C]OUIec:&d>?E[.EL+&\\4:2B<QPAQY&Ma
// ^+a=C=DcS:7_[/>fFAN6OES?5Xb1T2g5Y4FEQ<&>;86.e?38.VIgO>@#R9^QH=<[
// D>+=e&#FRgVA_U7#d>NX\d.-c3Wa\@(gVW>T+;+3/g@?&=P6F-;><HLH^Z/MLgND
// 2COO9b===45N#25,&]39V:;@b@5KY<@NO0X[M6&)=_[VcPX9_RXcKb?T]7F\\>>4
// #IW?BNWU98g9JX,1LW?0DG:X.7B/[-5eWK]RL6])U/7<L;L)Xgc\L;\a0BSX;=>7
// .9:I7<<1DQGE+Da?C.e;?[\=)H8)>>6&f=.S9<JgFP6X[O@>M&5MMZU\fJ>QfYPN
// bOTQF;F,0<ARP]P&0A,YVB-[Y05GcPH(&>_CSfaJ1BGf4B[-#&9ELZ[?60=&dCX/
// Q:AJ;cXYY.Ge<9C<(e+Ig/<>NBNJ>T0I[M6eR]fK)C=Q;8K?bB)cf,<6SH=>,F5e
// .8#aF@dB[8HWCU);SC=4<E<S?8Eb[g43eVMS?D0ZHDIN,\6IFf7aLb[Z1[=@,P^_
// c2SW@^9^9M.(=532RM90fE>N0T,KTHc3AE#[55)d)K7G85+18=8b9^:UHc1L0R].
// a+=Oe=,0?1W<GH^CH;R#X6H^Zc.2Q1(\S+VRV8U1C9ITd.PdLQM9/JR4]cS_R/](
// UOS&\E18NP?E/?R&K\=NB(dXH5,F.D,+/GBS51PPd+fb8_6LNa(Q@3[a4K)#)FPL
// 5ORQ>CLebW4CUL,E@\JPAd@7Y\W,X=]@4BCebd7ERU1(RDJ:QTHN,-0g28^H(-bE
// @@>0g:HPI#7JLS;3Rc^J0RR&g<acBd.f(QF>>[a/Z:^T&4B^ZKaS>P/\EUIdK3f\
// 162-DHeSe^UCX4S<c;;+G><If04AU=^=K32,.6<K/\/U?NOQ=IF/g[8-LR\gJ3-4
// :15=aTW&Oa4Hc9)D,bGX/6a1@M96Sd.DX:40TNLS:<;eV1_.[^)?ZORF+MFEQMaL
// da94FYADNb?77W:LF#^f]1(=,C04CG/#&#cN@f)X2Ba4OIXCM/eXB_5D1MFYM>R<
// [C<a&Zd?TT&0D7R9.:WeKTSUb7.#g1?SH?NAM)D=/;^=MDPW6/]@DN&75A)F+PO2
// bd\;KC?)NX8f[,T;W+g62P:eJB)<H8(9@4QI^BP&#8b0(bC8,SS=>R48A[6B_P=8
// QeE9GgJA.SfTaKN_Pd3203fd4N@X8a^08#a.@+Q?F6,4&#VWSa-Ie&aHY7&>e<E;
// _M=JA6--RB634fcZ7Q2,gRHY2C[7NXA4Q^D-,aKe\E-]G)VD[BQHJG(?ALL(\cUR
// Fb.J^gEgNL#)C:3dPTAcOISa)4)=LYT1E_b9QLH[@:HIeL@OT>DSF)^3U>8Z1FRF
// &RM-HHTZOH0c[Z+MC\]HeX.V+5XGHKD25Y)5A9DbLdW)M4.IVA_d^DYb8,#,f_K#
// f;JF=[ZIWT^6b,S@b-Z+5:>HB7S0OVP9HWQ<d/3Q.\fag094O-6MG-^K6FJ(f<P,
// .-fF-JJ,<49V.SO473J8NN998X#/AdaWNS+Z:/gcD;M&8BFKR>\c+Q)M_HF\XC&0
// dX9;/g;&9LZZaO@8CcU=^RSM)LU)Tf>^b]gdU94H/7M9&?_6QKX6b+\07b_W:4_L
// @dAV^afFbAU074Lg?_Z,b2,Q8K8Ib6QYT<=7C]Ha_P6-d9+OW)DPPebTIFC,+1dW
// ?VW?N;GVEb\g=X^YD2d;98,IGQC0A:)Rg-<]^W#?HOb,@V_c]@5E1(B7NAJ8I2cJ
// SQALfdI::G.:?1A.b3Pff79EDa=bYUc6/D]<_;OYbCY&e:0aUP5CgQ1)a8\::>61
// 56L+Ca)_1@dS7V-2^0X7+EQR<I-\cT4MIS@AcQ,:#M&#c0T,[A^0:>b80F9WK2[^
// 0W:7T&^??#K>+=R-af)0:LaObZ[VUNUQQ@>(ZV2&FN>;75O,EO-GFZ9IFd]\0_1F
// g(:45JSg,=_d2#8@I>X,bCI8BK1+F</EX[Vef8#NQWGE0IPf_@A/9)B[e9Q]d7Zd
// .+,:);[1BdC,bdBM\B5gJ8S#,8KGP\A>N()SO=,)2<8,NB-[_b#@?f.X1^bdX,1<
// W<QA43@_7IKcE?,]LeCHcVE/8c(5FGX#R10P?31&+f8A._GGXafJc[R5C@fbQS5^
// <OW.Ig(<4_/^-R(FP0M3JBaVDPF/R(ONE;=D49cY?=@E?4)>LS?Uc-5J-F=T]9?-
// Y_50O[O^(YU;_W&X=KU.PJZ=:K.2(^Oc=?S.TQ5664\#E1g,e=+I44OLeDP3N1QK
// <;.@B)6P\,CQ4Rb+45=44/?6@VUOaa66e2Idf+SV2W8#B72?56^:_cM1OVLT7;G]
// -U#\5gW;;2^aJ,+N#-[D+HWg;FD3&:ZRK9S+:RC1YM&/+;G:)RR?cdQg3G_I-S_(
// M6R@b\aK<ab5eP1TRg10:eZ>_Yg(:H6@Id5Nf+H?f5J&-.-:7DH/YA/2BO/+ff.K
// N0?<TSHa\Q^&GQJT8Qa_S\Z+e-K_3<:],EU,HBG7WW:0AC]^:6c&:,)O2^;a7;4J
// ,]Q&7=<X@/JN-J<TW=06cV9^=^9Z^:OV_VU1,3V<=f+H+KOK[^WOD,bfZ?0-dV+a
// +_47JHDR^XKV0C/591eOMB=&UMNH-:<e7Xg&f8+S\D2)NVLLU2@44-:C,+Ae<-TJ
// cNTg2URY>WTTfEQ(WMPFT?4KbF7R7L>73+2&U<Z+c+I/dEL;<XfRP,7(6@Y^\>#X
// 6dI;QZ\aJ4_V0df1(+L<b]g#PVRMKLYB<CFLR<1+I_F<+9\X#G2:0[>/B9E0Qd@.
// <cF/(P_f+LDMCCgQ?YX=DX6@Nf(f,4&d-d/2EeJQ-8T-@;MD2e<;8#S7VdWg1GeP
// eHd)82(ZOUO@FIY<Xd\?4dc]cG-9V6)bX-e148[DGaJ22B#TT,N-Bf./g+E8HgeG
// (]AZG3Z(S8G]S/fg8N&R4.7N[\Ne>\R[B#TYN9J<H)aX-G(L=BfH=9G:K=+@=1,,
// 08AFDaXb<M9Rf\MMf_D1K1PG?FPRF3H^=:7,[SMSARb;#Pfa71WEQX8,[VG&Y8-2
// W^R#@;PTT.3R&9SYPY,L1LG7\D[&?OCJJ.RcVIB<bEDKJVTHFbW172721\TdEO-8
// ^a.?caJMBVPBG_9aK]gT()I[6@ML<^Kf1+cQ#P5=V=7[fg(GV-.TP,5R43_2OJF=
// MM:F&6YDE0=H#0>Y@KCHeYR/-40[=ge]\\M=PZ_<TAS];8JVWb/a#Y?[QS#W,e[H
// Mab5^+f,P]9C<6gg9>)P7:gX/C^Q4?CL,X5P5WFNQDXUCC5KG]F/CAHY.](3:]K[
// QR&?He>3JRGDORA4[67&VR0\D5@20[R&H-a3?Z=ATP4R3-W6cAK3Fa0G?I72>eP+
// @dKFBUe[L:&YO^>WL02?_^eYf@I3?^cA8-e/ZeQ@G8CQPgFCYH+-]B7HN9\-4aO+
// @JdO7:f+@W^LdC\fUJ;0LO#cfOg<Y,>&.Pg)Z:=9X:_K(@a0JN)b>GKV1QH5c1(H
// c<DI8^1:FLW07g;>IQX0ZgN17DK]Fd([G9.d7VZ8BO5.;L+==FZ^bPWg^=-W0DF2
// F_>eQAY2R3D7<W/._FOC,e#W#aTIGIW>+BSEY_XAD?)&-7-<>KR]G#EEL)K;D9FC
// @f(B;Z-;2AG&9a>5f:SJ&(f3OU<RJZ[2a:@LTR\eAJ_/fa<]2Sd<&E1d_7>44820
// 9<DYC6?^3d34/Sb+MS=SS/B:&\NR>H0;/Q,P,((^CS.13FN.E(Td\a4PL_H0QQ&X
// Z^6We.A\SPgKQAHP7U9BH5Xc3\1J&];P6EOHA@Y?:gGQP+E7.:VZ<Z+@b\U_E[7D
// fMg?[gI2[9QBC#R7gb^V(#8#PW2P^Y#RW3cfI-2E(FXI7I9=gf^X<AUe.CI,Pa0M
// @-cZ=@M0>fY&2&6&AcN,=KC,(P#(eaYW0<_8I-O:&0(+a_Y<G>M.)4.=F5D^,WE\
// /-RNL++)d\YS>0I[-FIcIBOS0:07AR&U^IbG2IgP:?fdT3=FL-WbFg4Z59,Y\;>)
// b2/O#,GLegc30[QR<d,c1K?EbM+]6(;CJWgaRS[]begFU)F#aONXZ-<5:W4d@T[K
// 2?OW\cf3#WRT,6>F8]NXJJ]c41(+0T])=B4+)=?dX7Ie;^AECUARC#,^A(VR(2?/
// fg_<T(fOP/UFA/-c.P?^Nf4X&7:RC,S^RCAJ_e9W3[ZUQZR,G3UIW>8:TR[Q.aM^
// NX;+Z5>gF;f5+C4_10I0c&NV)FHgUQIbe^6?\3Q:WEMJH9QQ]cE/RXGWYKM>I6U3
// 9?;)b+688,#IgZ7e]XL:(-YAT_,<MJ^,6\gCeRJ@HQe)-c8C&,J,)_?H,dC<eVdP
// -f?L3S-73P&aS1_cS2_WT3OVdK=eEaX>@,=f0:)Tgcc2^8Z7G[U1@3:,5FUAZ(\S
// /6.<G&F(_(?EW;S^_32[P,6,^L=K8B_-)ME+&5H\EI=SA8PaTgP;aaJMW^K_@IB/
// SU]6U.9/OVS83_T.GeJP2#8ODZ@POO,D-2-I8MP@P44b9D?&#JBV::E9L)W1GSC#
// EHXf:K&5>WL-@BE)2DTN;+G0;]EQLBbdBCM>JV(ZC[@FKdH&3?VdY-_>#B04L(S+
// ]E)Q2/:@HAWFFXJBZ1+^[##@NAB?H-1\9?/+9QBf(X@0VYfJa]J,Pc-;O/VAK(a?
// YK&@VHT^#45]\#E525dE2L&Z7RKA[IDgb1?1_,2OJNKSIEU6?O^fIcSb1=PNO_-E
// 4W^K1-#>Td8L1GII6D@=KS]L8&UN1T@;,&SfcMX:F5cg:?9cBd)_]cUaeaOV/G<,
// 5AEA1JJD,.TR@J3f&:F;W^]=eMe-d:B>=US>dH9A>]G[&;FR.a3QU=7FZWN=3.=O
// U.SR&Qf]V\G0/I<?YO=b:D@2dZ3_]^HZP)/EA7K)49A,A2aZ@GZEA)(ALd@#dM=;
// E\/K8JXFAMTO:LNLe_Y@gL8d_8KdI[Cb^KbYdUgLAW]PEHQaT1,681\gCVWE:MNV
// :5F]FLX\\</7#ASId>G8WggHX;IHe6dc^J0G>g;C#=,[KC<79A?-PCM<33?R)XK@
// d\,.F0A.aKR3EgbB9V6>/B16&Qa,K,.F;2O>,@bY50[K];YeG0QM]9@#Y10P#[UO
// \5>31FK<e^I-^]PX2d3dB\^VZQC[&1g/:4cc:Nc_DQbD,<XS@_++Od16V6QDXE4<
// VA;(DII+MJY.AP&@,,_3I[K+V,B8_\/,)\F3d#9g=1R]g\Q7Jdc.M;16C=?;?CF(
// I#aN13Ob)TGUf))>BUS7Z]g++;&ZG7JaaeU[DHg.-4?ZKM+LeH1H(eaK8FDX]=VG
// f3g0FYY_L7;KNg@AI#=>adH8HFX0BJbKL9L7N0KNC\g?#1JD:C\L/,C.5\]RfH[a
// JDXN/PUd&)J3LgdXZ2D7AF]b0_S4bBIT\3;(I.TG]@]GA_]<TcB_52ddWa3=WT9H
// WS=VIcPI-)0MTA(Q<R7c#+6-#<UHNN^:76JYA&]V(c9_,\/)UUN6cS#H+Y@KZW2\
// ZU^X+)R_YE^4Za@Z;L;7)VN1a@>;XgG_dVgR26MNdMVPg@U&9TWFJ,FEZc1;:XTJ
// ,PJ@G3=R&^d);K]JR;0:KAd^H8cOWK<^b:c=g]a>e[(K,5XIC?/3R2F?4(0];]3W
// >K-X:,T2/fHPVFCD0PgBeL2SJ>[]:734TJGR5dgPA04H9\>I#NS>KD@06IO=63e@
// :KXX4QgW&_c3-?V@2,f<a3=9]SVUAPa\#/S-c:CZ@HZ7V.d&WHMT.:aT9-KMP,.1
// X0POC\LI9Z^-\C(EE6U0dPE0_R)+gN:F7fQ;+D:DN8[3>)6Yge50U+?4EQ#P@SQE
// 775A4f1V)J1/S2BCK1;f>\SS8Dd]e:DV-TPWY/0SLZ3f6<NLYX[5ZQ<+Id:18JS#
// )=5V^9W8bd9.#4H2ePEN=FY:NT<M54D-;9Ca[5fV9I44SRTG85BV+;TAVf@_FRUJ
// 69Be)g,1#EU(DRS[YMCA.QPO:D5^^GHTa2b5_C>:,YUVOUA7#B[TKN@HWC0KfAL4
// FfBBgCa5@.)1ST.R2>CJC,g?31Hg+N;NI?7P8Q2<P#Xa0?R.:X<-2(3eUR.)QMGT
// ?#]GTHRQQC[6.##[K0@cDd:9fd^#8QTT7AaFHSNF3eM.;64EU^A#QPL<EA8KY.K&
// g/a=_^?@VB-\YfSe:CbBH+^G)/DJX=8M&><[\]eG?M5P=6O7ZM)EC\Q3RUgEJ-9E
// ];U:,:/O&Y_.?C][A/;(J?S,0??FJD0L0LBc+;?(RI);2,f]A?cN&)DcED(;K[<Q
// PBK;84/LJ_CRPeZM@/=+C:3V0(NJZ>YYFGUgGPWPYF,4[g>S=eG/g9H/QN(G94\?
// ,+2_Y]?LSJ-2YL5CebI^Yc+(Z(UO4DaA<BXG0<TS@2LSCWTG:^LU:82;EdR;KNG2
// g@O^Xe^]G15_GP_HbA>M=,/>TXYKJGLW=c;b6<RXWH2EMbEWJVQB37@H\2Ua_-@/
// 1NG\UU)PU5547J<W2\(:)<edIdW<_3G6#I]+B[.cBOQMNOK+FBg8?4:F8]BSCO.c
// _S.3^YL+Z_HUL-SZ9Q<KEQ)>0eOS(@c=IH#_5K8YI?Q5GJC;ZG?:]WCfJK<[7?-U
// 6BF\V-.O)IYJPbN+ZeIVWQeP:C:WeFH3J2MJ6Je,5Tf=eGA/M&19Vd4g8Aa8eOaE
// 6@B\JY--Lb@H6e?Q[aO7,XYf>#GcH?N4bY&7)JC<FFJEPdeLVgcIQPfHL4)H)(1[
// =(dB7Y]dAe+EV@54/K3YQ5JRG)cY.C1IAD>NL_?5GCQ4GMVbBF[NMY-2fg./V^b0
// I-.1\+a+Q&MR6.&d3H^YfN-1Lb>D(SV[G9c9C;AaDC)5.cU2A=S68gEMa,]cJWK[
// _\&6)3H:MN5,LFV\S8eV>OO7B,UPf:a:6XR5f9IdH)_Z#8BGPQF1LKOJL41#W(6F
// R&&C4##IWHTd/b;?6[Hfg&<H;e6SE\4-3A9/>&B+:cX,Q@;eIUC]Dg1#3/5F:6PE
// Gd7J5Z#6bBPT@R=_bc>\4&1df7E0@Cb/Z9c#[[CC?JYZKC;_.BaD1\HTg&7KAU9V
// Ce(FB#dC4,#>62&#<CN)]ZdW:XgAO^N.7:^E/N1LN8J.8KW1edA-CFWD)WWJSK96
// /0bA\TCU#BL/b@?ULKOM;?C/V-+QYK_&=93fg-Y^I-E.:+7I8aY=@9F,J>:^fLFV
// VddFA\\Lb057dQ3&BDYZ/G3U?G.J36.f33,MO:C7P^6ME#LO]E9BN):+H1.7GH<M
// T)[<D1&YRPTG35^7Y8,86[2EUI#]SXg]<[])VBXQ1420?6A1E\>f(1OBC\aJ2_<;
// 2NcI=c6>B?8LLJM^G;OG2&4E+Z3/@,TS8eKEE/+:Tg[_,[9b#[8b?PN63,W5K&O-
// 3GB^0TV)YZdATU?T_BEQJCKT--.>DTZH\(M^/SL8>:\_5&KM19e6;M5bL9>abSHH
// 4>-)(+3#9DBZFLfIU&J9XCJ8]OTK;dF(S&,,OgV#W=bL:g]#)@+<O;Ef>F&FZ7gg
// 0[;DJgf[.E//\OCCG4Rg4Tb(RVV.R;&2:JLDVQ)5AI4-@R5#61#bA3]5>?e?WO(B
// RR->:aPXcd0Y+]0faVaHVULRY-S12Y8K[Z0DL1(()3<V3V,.8Z^1\]fY5_3fS@+2
// aI>DZ2..]O-fce5C\[f3=Z9)&)JEg+3L)b0Id[[.][[G)A5=@J]-S>-53YUAN]O9
// B+_FA.1,#50Pf/R&;29VWC0F5MW1QH:7@a6f74O,#ae<ba?dL<cRVdCLf#<>:/9[
// KYV>UAc_bJWR@8]4TT,><9Ng78PKQc=B(ZRFg[<F1>Wa0P]50#cS,6[M9W_e472.
// )9/J]bHaHaA@MT3f:GJTO9T=I2DcQe6R+/+\dMCF(VVZ\\14O:D/04(_a5f>\;a.
// )4>QHQ2794-TcWLFfVM8Z,1SYAL]V@H,W=W,Bef)(/LM:?Z)3/1^Q<6=DZ(f3X3E
// NX>J#.V?#gU&>PWHe75UMe(WM3DQ-;#?[EXQeM\Ag+Z2:6#Z-):-L=Z1C_MLYPQ_
// 3N@=@]Ib?T+E1A\6.29Z@a(J>dVV7B&U<bI+4If,IZZe]W,Xdf=<Na=M8Z(#]FC[
// WVC8KT+MJ7a8WaDYGgZ/VC>MY@NR9>V]BOJ)@eI<V;&YeQ:YA8V<:;&b]=5-K-G[
// Ae5<6?Ab,62@Z<?>?D8581J/LG1_37XMR7f:,8E-\YLReH=.7A+/)?3TLA2\B5LI
// Q&Y;JRE1:7&]^:ZLG)f2>a/_d(KHfCAf0Q+)KfT[,,8<:1Nf1A:?.;Y\WKc,ZCa=
// 48dCU()8YNWR)V;&-I/S9f?1^;^dDK,.G_9QTNV-f;+8(4;=W)DKOJ?=[ZQG14_U
// GF@,>K)3CE3C(F?19A_S?_cNU/(FTVN?+C&AQ5_GG-67P@d)&J^3+I5BO:DJGT2G
// ))ObI^&L0dA\/38NAbC(<AYW>bQAAEH<A1FEB0FdIGVK8UfX8R;EN(_#Q-0GAWV&
// MTFZ;7dV]VW:N;fK]ZB_:YYDaXQ2f=aO^LVJb/\ORa[ID;;[95]5dO\GfNJ0@WTL
// IA8b:G5^ULg_NB8MI0GKH.FSSeW7;\(VO&,CI9#75PYfg@(]KNZU@]WLB9([;4V:
// [\L@5A@B;^=98N<YT:U(-O@7gCE=P+cUd@.d7K^aT]IQ#:RT9G+\^b8)77PaIG@3
// /9N\?E<cMC]d\QU6\]WA8NgV&E+&MGe(;P[=?9-U<.F3g4&QVAADNMSbUS#C7-&7
// R5VLZ^7:H.C7;Ab2@KZ-H,:P^)G&H.dSIHDe.3Q?/(<NS)F[H9Q(]MR[P@WH:)CM
// E4^U\5/S]1XS5.+g2=,[.KTJ]#-:.Ge:J\0G78b4DB[OgZB(T9R+OA.XM<S?1H;a
// G+K#0#aVBVLaT^YUfKFKU/W:M9=6B82/N+@OM\-EZ@QZ=_H,9[STVI#B:+VaA0@Q
// T2]LJ_CNSA^]Kdgcc9#UA&.Y#-CQ5cgbPf_M#5,;M/DIY4)(0JS_E(749L=PeNX/
// 8J](8RGedSBK[=EPgf0\c+Lc=a.O4D6,EbC&d-PDOMe(P<PC886<.RcB4V>/LG9f
// K7WbT:D8^XDQZ.K/#Ae@&KV5OC3_(VJ,;YEf(;>123D43\=cY&\e\XJF:&gZ1aCI
// ]^]]K:IP[QU6c<04fIdX0a4Gg8SFHd-_)UZcf2b85V]B[g#=6O@>PF0+JS#1NF2.
// 7>3>=V2Z2F;Q=360OU9_)4=43;JI@4cEZ(-R;J&<L4N>[\bYB,F&D,I&=H?bg>PK
// J4C1#],-aTaWVX<NKT;cQ_0RG.?dL-dRe5F@cNMU6<&>b=b#+,9eI<XIP8]M3P9H
// OB;239FcQD9F4GUJNe2Y#X75TCEe6:1JVL85+bgf-Q41Q>AXL)>ac,^fZ=fde<+C
// \&JY\4C)X9PP_2>0[?W)9(ZW07?J@FN16PIA;7Q1fb]YHgYF>YTc]<g+fFaJOODb
// JG344Ac_#;;6g3#UNX7<H\;K&+MX;_[Tg/1_E8RZ)fL?[T^0^TMBYAH>&F[5:/b\
// W)M^.b_JQ=:Wg[J)(X^E4^76(daV_7[;SQEeNV2agP/BJZ&MP-bFbN./[bKVeIBH
// R,S.?0+GO6E[d>=<>\(NU-&FcG>[f<QeQCEFgb&SQQ&:\3VJ6X62O:a@]gB5VT2?
// B,#POcWKG?<X&[_L,D:.501aO(AXAX1\Yf?<_B3,/?B2?Xd;385[)E:UQ0>0X(Qc
// b-/2fSO=9VF9JAX0:?-3_==E,YcU<bV+=gH_VGTPC661@S9?-U1;_EF,(GKN=#Sf
// 9K=X(NW-9^.Bc]#2f&>:3THNK]_:3HSI)WFW[J&]XGH#8GP+UNA?ML2c1A]fJ8Cg
// R>?&\#f0#e)ENQ4Z=&)YXECb#;eOdRFbP-W=bC+gFYNT/<]D9aA@VZIg+J4G6S/.
// <&(>cKUN&0?S.C3.UP0J\XdVgag-D2.N0#W=Q&R(+-KUUT:SULTVN+eKJ?,5=)R<
// 9QbPP5CJCS<Z&;B&T@P^5)#C)>QdBC_Y]bB4H85aS3I5_6<^)ER<S?&7W/+V+c-A
// 9MK14?G-cQBZXDYMF.dbb0R?+e^Z\A95#@5ASWB8cO5cLdK2Jd#MaeN(K.1@f?Qb
// \JBFKaPbFII5@YE3]Zcg]BV/K=RS)3ZX1O@OA3Y2A..6@JN.KQ0@ZAHE9WBR><[T
// 0)?/a4RSB+>9H_JKV-C-2D&BQ4@_/?P^[H^@>;IL,4N#g^fdS-1a_cJ9A;bUf6@B
// T;V(S;LG-W(_HGM/,\UQ4BWEef4a:C]49NQ)UcLc+NAfdW3?9X1:</aECHR@L8@N
// GVIXRdeZB(gG)0SM3(T#,4eUF=I?#2RH@O8M-[1H1RBP4U7aQW#@IS.FSH=Y>,Wd
// =/aYEXXXdFcNRb4]\O):>5@(FXKU/I:W::R_b_[BAGVA#W1[-[?^(0\7TKZ;g&5N
// 3WFEb9gOe7.I1dH_4Dd809:)A-@5M.JD0D^f7)?H9G/dU#Q)[ZA>S+:YT]1^VHgY
// B(T/>QCE]BG2;;#>6XQa#UE=I5gTVAEB&T<b3GT#NE/dT);TK#MJ(@A)(BR?[EEH
// AQYD&=eX;f<FeaN;>LaJcYc&)[eaH\NT49?VJW7Gbb+B[D+KA8<c_X>Y.9de>7O8
// R?^=BFT^Zf?R?;8-=<9]G4=4EK#Q+,4#UXBG/eXEJ.Mgb_DQ52Y+KMJ.,WNB>NDI
// )BP5=BGX/S^OGbJV1(.EUB9<fDCc-gDg-[RX9^a1+[I_1,OB,M@]XUYGBMJFV7@:
// 2DW^^3)e.<I;c(NBg_?_7RYXV,RYRMRJUCVT-7=BA4F#HL>9S0HF,_IN/PTNU)A2
// M.C95SE2#2V\X5?4cTgJb9^M6P+JRGWfY,W40/FH#FJY5b6Q(+I@^F?A?b:#e)?=
// FABgbfg-aIM6P@V=bX>ZT@a:b5^;-4;(gJDfcS7E_>.U+37YPaL:U#7(P5@+Q_2@
// W2Xd9.)[EGSb53?_]COAN=;e4-aQ,JFfd<\D.\I?F\H<;KBg\61H(W&#Bb+[8SQc
// [NX6.0cFd<ML;e#645dVT,R23#:(XP]I<L94MbQ^I#b-()g]ZF0JY)fDJ1e@)A^1
// ?P_83(\WP_4.YU<_&L.JK\GI]8F<D)V@_P57F(0(GeT/?[&T[ML7HJ;XC?:K:VTH
// /(H+9+&O>K/?RY>eW=K517.W_0eG)ade:BX21NB,&..b,/1LA^RV_eHCVFHQPM3#
// &Bf1WH?cfd1#c4aGK]_GSMJGM1##QdX.52>SPNFG+P7<FW&YC<TG)b0H(GVeV)IU
// 5[(8G)4c:?<b,;J>ZAL888b-1QE.D@K&O-)[;;RD(#W98N@U5J2TD04RW,WRSW:M
// U4(ZR_b](e^<[YF_;_@)+#:KUC6:E-IO-ZBJfAP>Wffg;80YKVA2+D[62U9SA9-.
// 5cEII?N9>cS+Q+U)gBc&:VQP:,6>QLZR6Y\&C4;5eUf#?25W+5+@;.Q.KMW:fN:c
// ?H8Z&HH8ga<H5;Y]<MQg;0b5ZYTC\;^7HJ)?[E61XO@=]NX5DS^^Z&-SAYL:DW65
// P\cWUC0d3UAPW<G65f##&0W:ESd>(3LH]e#,44PIY-8EcGXTIH,GV-K\?]?.#33<
// b5H^Sd7>A44>9YM5R@;0:ISA2\Zd.;PJV_.@_UTI&\+F_;>+<@BOAaTX#2<9)40&
// aXIR7=Q_\@SPDc^]/a1DH(J\7)@^=cQfPbRJW)7:JM5S;)C]gP?AVM).PED^XW._
// [:W1ObAWKU4bUQ7N6g2D>+3;U<I1TEC[GY.]cSY5=e(?;PVFfF&#e/cNB-G?2[N-
// A(+Z?_NK\cMa7_80)VSY3EEB6?)fUf+>@=[Lb),,c83]IcWUHEEZ_M>:&,K81+&4
// K4JEfMI6@OUB+<99K6dFd>g.d;V=-LI_WP.58_=QM6KP,YYB/W0HbY&e1()JZROH
// g3636TQa-6QX#>fS6RG@.UQHB1.H9;HX#C#LaYb^#ed]Q&V060cX9aE-,/eaDW[R
// ,4=9RU-_N=b\4)R/d/1ePB-Z4Z<U5BLFX-4+Z^b(A=1W=.9Oad\.#cJQW\=5#,)2
// g4<M/=G-dV__6eQ,PKEP1O9(;Dgb2H=Qc&Ed,UV__W?D1DWT0A1^PM3HS/aU9U=X
// KgNdDTAdUW9.Ed\96aYTY(ca?V>ZTEY:^_;e^f=@c3)e^YBdFVMTb&P\aPbU_RG-
// I5J=[H-d.M1=I^8g6<4KD6S7A_ZL03P@)F@;cIV,#c2J[C)E>6Yg#Fg]2EaUIUAc
// 1;KT7DLW]+c5e/a^c=,L(?3[JD,8,9/,4.aZ79-aZeB[/0W>[-A=G8QYTM=V@R1R
// Z6GUF^QLJJd/X+A7O1UCIBT=T[1O]DaBKNR>LLJCc?&=GPXB/YFE1=GeQ-QVF(-g
// \.2)3K/R)59NF_3>4db0RUCEUac)1[45a=d3B<MS(CdT+F5I4G.3Y,9D2#5Q0@fW
// ME]_I_XP2c];-aXVKI9_RH6W?M,EI_3MNE3T?/&6#^B[A.\bIKD_GBdX4X-cV3d#
// ?ZIAOE\c+Y5]M;Kc?<BK=3e_/P^)a-;C:4::=f8A3[DW@c:Pf<\3&E\ddO-.[2a\
// 5VLEP)F&aRM.;;c+Q#eNXY+I3E(ZZ[+1Z)@VTRd#.g)-b71(MI-YLBRLLE4U9P.N
// FJ&1ULK8;G2BcSTc+[3A7fK)5E/2HMFb@SU_f8#X7Z[6LXY7E33D;BOcc/Sf9,9/
// /N6W>&7@\S)G[_?9.-&12Hd7@[,_DOX9GcVN2YOP^?6fcL,#?SKV^&<95Ld(Q.S^
// bS8=d^8)P3HV/E;g7J+\G>M6VSg6SAe4OgXJX&UK.<HJXN;1Y=#.Uc/=P>,.SYbb
// OHKECc;e_UA>HFEFe6,=2(7D#A7OH1=c4eG=&1C\#ebWSBB?TG6T2X[2-RDC+8SB
// A_&4R+g^>),0+B7fH7L?(T)K74\dZIWJWfZIIUQSAV;MRfF=Dbg4O((;Ia<>a3<\
// E;+&:>-D1ZdMY(H^aIIU&]P_NEY1+B(gD;>=7,_SDVOR4QXPW??bA<:+K:]#dEGO
// .OHTgC4)daD(f-M-dfN0SYHV<Jb=16#/[1RLL/5?WGZI8GM<K4Eb=EQe9g2NQY:2
// b<H)@@ZcMX0F>5Nc-Zb>b]\QH474cD.[,,WLUX0:SZS07>9H_GZ7U7c_]S2YaKOO
// cZAONUN=fCa0RHD/O;6Q<g>^P,dD.f@Y\L3?(=ce,H;f(Ob(@7@ND^Xac\Zf+0MZ
// RTUH)JT[SN.5RW_]TQF7eWR=#IIMDJ^C>2a:J\AN123?AV++H^(]&908WaNZH9Vd
// C^CIG;:V7#b2C)-g916=EW>9@ACe;_f)c&DG&gR\a_ZE0CPA[0G@XYLfHR,1,TaB
// N,a>ccM-USHEaX4E/b8g+J3E&39ac@^B:TX/X4M.RaNeI[?6/1^<>#0;H^B>16]T
// d(3QZ:8^=?]fI,4MCW=\^NN3O\RQC^ZbMK78OM.TX:IeG;](4JBY(?#7\T9=c<@V
// ]FbAWb>1.UUMU0cZDg;MO#/6N;N)>e53@.0bQOOfT-/F^41TFNYMU,]#Q.>+g40T
// 7B.eO=>JOAf+\],eE0[6TbHbYDNN::\(d^>dN<2&=FM]PMJ^b?UJ]:;@Ed@2_Y>\
// <P::0a6_6?O4@2Y>F7Q\BccfR#=_S.6O.aa4)/dV:H+ec>0&25P:7Ff4L[KMWP1[
// W>gN?[GF>+\-(/)BOXRC2(RSA&CaMJ=DfW@<@^LN(fPX1=D+G_=X<g)VZ&1a.&#P
// @Mf,B.-g,Cd^K[O/A@c<E2cR3WXVR[\&U4X&3+ggF:WJU+5M;<\GPc4fYF.Td,AF
// /ae0209@7Z_@BIFd5O4Fg=-fg:LZABOPFE@CYO)F/AL8D7<.)b[&4B8T@/??N/?D
// cAI=ZbU/-Ic&8C_TWc3D9EN5);8HI.=2<4P<[&e72JC>HD8)(W]TfSQ>OV1<PWV<
// -,=O4bONeB<<G/])Jd5[6WU187+#SBZZR@Jg.\<FR7#F<T3IV5Q)P[<YG#GX&67[
// G&@,<EQ&0f7YGfdBbgf@1C2S@06eJN/R&<,UN\-.9c&>_5O4c=Y.G:R7UL.I@/cf
// ^A1#8[Y:@+G?I0/U^=Pd5^YLSaEN^,OAe;9Z3I3&?#(cKSWX^0F;;3RO0K6^e)SF
// -:T/_R4)H#[8ZZ=DNEQEM5=g];U;f)EV:b00(8\]BYfH#ffI9PD5IKPFO/,b,F>)
// =>7g\gfIc+0;=2\^+#(g1B7=.X/L;[Ufg3Y454c]YU;4#a/^U014[WM<T&cJ\J8N
// W(H/WS44/1feX7Je0KMG#NZ:?ODN;f:\T0F6RS,DQ,]EZScbC6V+BFH4^X&0+_YT
// EA_G8UVF:=LA04P_KOBa#aDT(<4XWK+W.b(+7DX<-?GWgcQ^BQP6RMS:^]E#T9S9
// &>TAb15-?<[F[<SKf-Q8.Ge@\;QE-S7c9b=f_WSN#\[cL1<G.-AeRP,VV7BcO68F
// 6XG#DdY<5\@4eRIY43[?dGbdI+]ML8>U)[ILUe&(QZ@S]BI5:XX_UaD7[)BT#H=W
// 0\/4UcU:V:(deK(ffe<8_H:GQ@G1\?H.E(_E.RS]1VXUba\8KQF[f&4^_6@O-=D8
// &7@#<##SR]4MG_Y&T(>1-Q#V5=(KUSK?b_c:f</cRF0-(B:f=-UC<X2N7ZGD>&d:
// A;K7Y6NBg3I0<Qg,8#W8CF8Tb=MPTVV9TYc@^[K8G73^L[f633<45.D[GZ0A]KPg
// J_YQQ3X=bU+EJ;c5Vc&1DbDYF?&26P.)U+QLF:Z]+6;/=7L9OCN@&>T<@<P<D>1D
// _gIOU90=73^XI,\Ge0eN?8aI^c&XfQ=3BP847e\A++?-GLc67:N4SK9Y-:ed:4>2
// <X>OCK79GZ#bRJ<22e+GbZWR4QIEaOeB8gb^;EUK,J4RWe+:J<MLNg1R_]a=)+4M
// 3TKe/KV89(X^+9,833@W4e6d]3_H6_A_EdFEePPc_PCf^#VJT:eV?>/9EPPEJUH=
// .B6,_??W@MR/B5VDR4_OM_3V&HW_FG1ab\Y,15IYCGHC5,RP)e@-2bEXL\bKBWDT
// [<a(]_@3_?bG7TBPOd/,Z\_2R=1A3,MF/;Bfe56Wc8V1K[=)L9<QZf#,P,/7#846
// [3,84#ceRLP?Vea2ZgQO>,4fJeU,a>)24ScDX=0P2EV^^2dIN8c,9>9G6,X#HOO4
// [P(A\IbYI@06TKIbO9?H\-Jg.]&0DEKW[;E8;1Ka:_J&eaTOB?-?R\C+.<-DDf;X
// )-=ZD-FF]Cb<VI((M_cKAXIRAf2D]AaN#/6=/8=<=Qa^aE,aBV#^>Xc@HK7DYXKO
// YWX_=3?6&6D#GE>K)/GFb]U&UAHW_9_Ba/;(<=JIg<E-)6_J2D(0:>A<HL&NPf(&
// 0AT0\4;-.NLI)T#D5,Yf]HCWO,C<cFg;OZbBOaVf7?PI?I;P/#UHZa_^-GeHZ=94
// WO,+3LVDRZWV>LW.+>8>:>;)/fP[/CB[RVe1XB,^]QCT=QHQ.K&=2MgS6Ke=0NEE
// EaIM5eJ3aV8L;NK9/E=ER&VHA2@&gEJ1?E2WX9cO)>+\#WKV\#[TBWOY34T^KM-8
// RSF#gd=9)^1]+H4\;9Jc?5X_cP2,1]D4Q00IZ->)_e[a8FJ.7P3#15>234YI6D\A
// Wa=)5/,F;YN2G81N#Y3173)#R:YGM?F>aaO&6)(f]\FCE#PC1[]eaFG&N#c?+>0/
// WNCd>0L76E4RJ&V;EO8BB_#@[TE_<c&^NJ?/3JZ3UX?E=FFSJ(P]#)P]_DLG9(Z]
// @L:FY3WBUC?;1<FYGJ(8B8a#Oa_(.=Nd+);<eF(@;-a^#@-OfF+-W)O6TZ/,^Z-L
// N_IGU/DI#&XN:Pa@^BBbSMDSXeKD@TBg7=FIU=>@5XQfe9K+X4N5.;,,(6dU=AU4
// ]NUaM(53bY0-POPW+>:d1?#<Zb2fMBOT3_a9g5]bKSX<16#R>XR@+B3GKa[S=4+a
// gL#VS=dfR/a^/DB)DZ^0J>D:_T,S<T]LH:]0UDd.F/KT-&NG0^LH5bBGBd4)J/WE
// >QW/ZaQTCIf\,bWCNJ;Og5AX:(T>#7].<RCG8J8?<WD<GgX[LK;BYf^N?d#;?NN2
// .Ebf.UeZSWaZIUeDIggDQfF0YH\N5OYS)+dP]eBY@5M?A43_X5K04QJ,;>YR1_&#
// (L-TJ57c_1VV6cK0)@P:4LV_2^62eY+QS]Ka_fX_<?3/g)=e,?e<A51YM/,W\B\G
// g[8[DC[@L4@>6Q>TJ_2c/4]5E;OYCOP=OOU/P/e)QEW+2M0gc8&UZ81Rc^:4O]c]
// J[L?bL(#9M@B=LE-DL@N[5gNfF:E?8AE(HW]0[-4D)-M+J&9O1H9db[\Y)[#H[T9
// KZGORQ.CLDED;II<+IE6??ZTPCZLI7L,^7g/cR#bN#4Q44g[:a14eb.Y)B[B?5<O
// E8\#0CgO=>IfX4]D>g&HfM:Q&BH@MNgVW/Q7\.c)9YFC[AM6RUD>]]G/SK>(LA&G
// Cb=.A@GQ/+ICHMMJ_2,SV@-SB)Q8LFMH8Z)>X:GCc[f4CcV+2)d:>MA2Efd4Oe64
// K1QQ.LF#fBT04A2R6@ZC3bSbJ5-a]bWC@(G<FM:AMKc)8WCCS)Vb)Y-?TdI=HaNB
// 5BJP.:?d==F;N\>?d[IFO4<F?gVg/8\+<cO&b_<_6P95Ja3gcMO50[bZ/?[=R=g-
// 1caC@>2Hc<S/B9G#\82N3P8)13gb][UBENaDa-+LF62<-(O>.,_RfX&0<BMSe>[e
// T63H@KM)7)04I(R/T>FT=NJ-FKO_U4ZIeO7,NdAI/GJ]R[I&VY1MKVW@=EN?4^@3
// I=T]dUHQF(TP<\]2@#8(IgP,4[]?PKES^E6Xa56DaGf-OIC82f^f,)3fK8/Z@L-a
// 6Og_NM4#UU?e7I,gcIV+.W36+cb&>:d>)\CUYbL,;[>XHd=>e><N.?,[34&PNY_G
// LU+b3W5+D.,9[Gb@NZ-OS,;,?Ub7>(]e1]7SULeg=.ROANfa.Z11OGe+)27-SBK#
// -\bMWN1E0MTe,\/LR]6,S]+M#^I1b4[C_PJ)J5,L?[ce^HQFL4,WX+5fV5L-=L.F
// 38H(&_,&A-(Za,H128Tb]]C8=2/<+?CO,Z-O=eQLW>;Rd#B-/C?:b:Tg1[;T(8K4
// _/UdC0P^AH.>gS[5K(MMcT<I+5/CPDN8GH5B6]Q.Z7TM8RcL+J101#43Y[RX(ccB
// #&>,BA0:=\+AfX5:)Y2#C(FL2FR,.M+d\ZRO14C@IgR=KP+;1>)aLO[V=:&9OFYZ
// 39B\4G(eI8)=Vg<S5@DdH)Q[P.(]Y8=.Fe6Y:N^L>.;X(\W2[=/T6dD^a=)cgIRH
// ?=)G@-O,#[5<IW,>E:\f6/N?@UPLN#J9_gSdDUg#Af[>0/;/>ZRI@5J#MdBV)CcW
// C/B(N>0B)0BJ@LD^dK>[S#P+F9/c09A:@:-W^ZP(ORQV/IUD^+&,I\T?aG^aE0PY
// C>eW0-:dZ[SSQ]f-1E2=HI:-//^O/PcDH#)?RM7H;04\VV74LfRd_=J@O6,U0EM_
// 8J&(+-7XW4@/WMFMDF2>ZQU3SFI+^@5Y7<2-[VP)Z\-+:c5eORBH].AO]I:(<d#-
// X.LdQ<[LY=&gW;Ed1^>Nc6bCT]JTb7FJYQLIaHNe[[&-@V_Yb74(K6?Gbf6=g3Ha
// L+BcGQAd(-W(0,-ZQ&<.b/6>02SRcR=g^_f<V,)=[cKK80,;RR3(FNR;/+Z4&B+6
// [RC1LC2Y0g,8I=T=?(UEZ?S789YW_+GA]Le),,A45CcIR0ZW(5/+L_WeIf9>IET7
// W@c@MeI(a0(g,\bO]Y\Rd]\H4MR+E+=b00=JUP.[W2W)g(d48QRBFTZ_e(Q(1GeJ
// Y?g(8)dU7^(TWZ9DW(a9,+VN6@;RO/gIJ@bgFNS_5)E/KD3G#d-SJ\K2JHDXgH0C
// ;b?fYK26,g(FS0a68/X_Z3_Yb++8b)+5]c>^GGTQBR7O&c6G&CY33BK@_We-RVCO
// gHBGeC:N4P#.<U(6[,Y7f[fKU;/bGHE4+>a5eK])V1O2GO-#QB@YR@T-\D#BFf4a
// e;=I0?=bd_c_9RQ#@)+3>d2f?4\,f.f)[aG3P:89IY<S.,LT+1cW>e]2e)PG,I>/
// .[9Z/MUUId]CRFLDMS=G9=&<bYa&+;U3#Q.R[afe>N&O\.=c<BHcPg=T/FQ5)c\N
// ;#<<Vg\7eS_]A^#84&64J<VA5bf7O^[TGUHSEI7Jb.@/L,;eM[-@,<KG/_[,<X(L
// NGL=c>D,G66SDJ5OMB38Xe.fea[;>Q=ZCE2NJJ^3OceWKATV((f8(,QcSa9PL#IB
// eS@RQ5\(G<#R\8\F(\JZ]d2dO#eHFI<HZWfX,:>OeE4gd,8:>]O]UA&-FDW=V+eI
// M2T=_48CP](Z_/E(4.3L?R1TZBJS>P9#F81/_^E9]b=^OP(DBYg5I@&53YQ41UQg
// Z6YJC1cF?7H_C[2&UXBPBZSd.C)D77=4]a=41c;4T&HA-&?9KUVM@15^X:OFdI3.
// S89IA:5^dE:c8.bMbU>;4d<#AFQ](6B^][2\PI93H+cEZ?[C<RKeU7edV8N&&>DB
// a99^e9M1RNG89^6#BXT/QOEUO#@dOQQP9g=[><SfYNZOWHOP4^<JMX[.D.J(HfQb
// ZUFXL)bE645a3V=dR2Y-eQSZ#=1^DAA3:PTT)DG>8FZ#D(Ngd2a;G>^8,W-=@A@W
// D8@_GVQF:+Q&W\/@XP>,KR5K;18=#A#;C)\8.CcPQe(:[gE2[_gD60If1,;X2Td>
// =J2;-bG6V)bXTSG_@>Z#95_7:F.((NcJ9?J:^6M6M_DL?(]&9+#I7K/D)DcS/3dY
// +4)F^D,:<\+)1BY^-,HV>\NTG7H>8<;H,//&aaVCWbFcHcGb4I38DO^A.&QUdUCM
// KMAN[,7@eRgXX#1W2.2C@N97WU3>.bedAJ^S0[\VC4K<DBe,@\-[X(7.cH[+M]^X
// J_AeHIKc9>F4V_-.XFXHSE?&4^S+=ZV6W<HW:<IXG&1+5-46b+NW4DQfIaa[MPRd
// eT8_UR8?V15UTKE)RfYgC<]XC.:.aN([J#=g&.Z@A@e_5\a__D\D<TfCYQ\R\47Z
// ,>c@E_Qe<WDa@]GY?&LA_0G98^)Ddg_V^[WbR]7GcgD1aY2F&RTfH91#&C;._\:g
// dS#R.Ob>G5._7-8UHQHXdQ\,^63^S0-L?G)eV+?ZAY42agSED&JG=O7.DKKI#f&d
// 41H)XG?L42L6@G/])A1J4b>XOV]=g@E^<PB4;^=65+NUZ5CVIJ#]PVLFA?N/K)Yg
// --^JBR-#I)c(@)=/U/51,;E6/GZ/[1WFg>KH5G7?P^W\ZKEMb<\/T.g>)TS.?R_c
// B(_/06F:b+fY+bWNR636JWg_KaQ?);FS3_3_EGYP1PZ^7acb6\=(_1@c7R67<M?E
// E[5VV3<M@Hb_G14J6Y6)K4OF<VccH0AaAK7P5QCW,XDSA,DLXCYU5?Q.7OH?-9+1
// )gXCgE<^YFNYWf@3d+a+/J)MWKS311D_Rg3[1[;Y,B?5BV34]<X<=DNR,LX-M@1T
// P#\ca-5Y/_QfA,-;M&+FLbU=2TEBY0Y:=5=gSXZ-RD>HgM:KNbdKEP9><UAY,IF9
// &=R)<ZIfGRe_UR\Q_3DaXJc.<&9#=3H=V:I/_^K:D9D1NIJf,,B\XSTcI;7S^HU;
// URV<Y90M4JS:8?6?=)O=^aeaOQ,+3-,RUd.B@P[c0[.X#U?YZP#Y>2F@LW7L2F-D
// L/4OEec?g?BFL=bULU:6>-f4W=IPg7#;+IG4[:71XC^]a]V2RC/a\F<Y]T3FD:cd
// H<R=6R;cH[91=0BVQe:9NATHG?a]H(bNL<=7PbD#+1_XJXY4]e862BcVEZBTS>XA
// ?-N5QT#eg2AK/F=Z=K,gV@dU8N=XJ_2a_#L#Ab4.Z3Wg,c2;Pa[fH>ONb]>gPGO/
// 7M^MS6CaQIg]PRZHN6:SUXD.H3/\8,IcQLHFFB<N)QBP3g[BAC5+Zc@5#T:2.Y3\
// CQG.60N62];RLAR.[AU=,H#7&K4Eg8P_^EGE;7BC.W^/Mgeb+5N\&5-(+9gYYfVV
// 9QdVIB&B@XDW:D#E4U.PJXVbVgYM+#aZF_U9^PIPE-&b2V3+_cSKY\fL<<aZbgI8
// 8DVB0FOAUc]M7>U_>Fd#BRB)fb9a0,H=V()B1MJ&LN@RWMDYFMTU+YIg7M^@e>(@
// N7^;&I-3P#Id,3g<.U,cW;D#/d6O>G_e4/-XCH);I&T]N+[fLD(<E@LT02<84^8G
// _D12_\7,)?&4[]JDFEgOT=0XY#C/:PZ1JO6+L4=H/&M1dJXL,+]&X[TK;Z5dY^E=
// R4_NgGKRC5(?9cP,ICfA-NBgN4.&e]1;D]1<T7M<3fI^WdRL8B^M50U5_#,#Xe8;
// B+UJO>.MQ&R/59J3U=K#bW(H.M9^ffUeaGJT8=Y)L:<2aRBWVPK=0&M<L?&EFV+[
// 4@(KI)]SeG;NBJNJcXXO6X9(;e8b777=J[]7>Q><9TTcHH\fgNN0FK9F.H(WIT9e
// 6(;MUgTF3/9HGd]LUg6WH.\+bLZQ^<V9/GC[T\P0+9a145^=;T^dLD@eB2b&YUg-
// cf9]MbX>^ZHS\/:@I#bWD?5?_P#PMdDF#SMR/R;5a>E/P5UNPUWQb(9S.d8OE+U[
// 3>MNC@Q-KWP-,Y\E69>dJ&U?PQ;#Z=&=cC(K)_D3QLLO39QCP&BGTY<;SgA-]HEW
// XddVgGa&#TCE7-(XDe799JKf8F2]e7-E8RM3K5F<2<^04Ka@N>/e0Y\2T+/gaP>_
// LC:c:aeS2MO8?#9BO6WJHB#JbRdZ1W7N9BR>eCT7NMe>BYHZZ+;CbK)>\QM+_)c\
// 4:&:)==D7<:WcJ?1AD7c+8N;1WZeY1Ue0<gNVLMU/)X:ET_NC.-5@OA75Yb4H0G;
// \7N65EUe4S?^Za7[H>6<gXJ-,YSe033D.c1R_)G4OFR462O6>R]c[-_)I041aQQ0
// ._(Z\F^S<_c,c8XID[7]R&>9TE0BIeKWO#DII9H2]DffTVPY/L-,QNEMI)^O[M7#
// ,T/?H^4.9=;]##La0fCTQcE+IH8Y3GLKR#(6-75K^<NQK,#7CS+EeVF1T_INNbJ1
// .&4,Zc+dVZ]ECK?_QbaTQF,H&[_-OAG_RNIV)&SJXLZLf&#=gK#1;O5<UU1DdS=b
// LMEH0IA7R?Ce77,0EWAI\EgNE6cNSSE[&L?#c3IYcBGIIXARCOYcXK_R3\(AAc/G
// @gb.fF?G;/=.Q/)#/ZU:1\KFeO[RfO[F4MW26YLCK9XYH-1<fS+LM^bLTBc;dD:/
// g/^^V+:P&Q\]/T2&/dQTMUQYE-QKILCCC+JT0AW&YbH_E,JXNV/\dH1NK2V-TOOe
// ;[H+ce(0[aL7O;.VX?7(3)dI)dW/3I+cJegGQ[e?&<<=3OK+ccGPAL/(MU41JV@D
// Ob/.^eQ+SS#U1@TF?PRc-Gg?V,DX=06CB>@/\;36Z1/C:L1/7e5RF]Ra]2^DA_K_
// 670?D=O#[,Ea1d.U9>Y-<[P(DZXe64cX);fC:@2+6d\O.DLWQd<658UCgZfX>K^b
// ^+:8[(&NU1Za1580=bTDf,3S)>8,//O>=b0)O&#?GJSa6M<^^B0J5Tg<0<K3_\aS
// @XD.,NTTPNA249[AY3OB#;e#IU)J.d7J&L:.]M?,[#J_J4])3,(VS5H_MK>N3371
// MA20)@gZ^HCGf:D(&F6eaZL[JQaU\9Z-W9TdKd)?9XXeg5>[-0g=UK[&IU#K8bG<
// 6<K7&=:])NRLQT]7g43\13fEP5BLZ[ff/(fAeYdUAR,[_eUaR=61[U):g:[EXN.b
// M8aAX.4fBCdIF0D/O0I)CQ]1ZI=)f0V+T_P9)(S^C[SW7fF>B^:\2O5]N8dTDg.f
// 8X;+b&Z20V0eN+S\OTJ/&K<>PHEK3^N.A6#f=P/);+b9.[eOMY@4:<6[:BE0=:6E
// OEe/Y;JELdL@^.4474FbYAAC<:f:JN9J#-//?;1\\_--<Y@B?-HD.#N/2AHQM8\.
// f3(>DBS1?D]->cB_V,-&^CcJU/BgX56bG)?0Q:1CS[?0(?\Ff)+\@aOQLQc=?9HK
// \Xc.T[6IYaMU+L+D)N[><ME,gR+J4F6)-Q,WR]0I.3JAMV0C12Q;gYZ1?GNI)EEe
// WdS]5>1SEYW-e&5c#K_<QV#BU<P9Yd-5-,A(?6]<0^//M=RFd6N_b\0/[<8Z&LY(
// #.ZGO8#;U44eRE+/d:-f^Z^5Tg.OXWgPX8/EH,I2N6[-YHb/[Y-_(WE]g0f4;S_-
// VW;;T#7P#8[]8Le7L\5BS.8UP8(IKG[(WNcEW<IB5_b42Eg4eW2+PA@O^)]caTaK
// Y@gec)FEVSC4<,e;ND)E+A-6(6T;f_?B23KXAb0@4dW8fRQ98YBEYEP76.FPe1Nf
// Zg3)9VbPD)]_YdRcO/>g3cg[))50M7bQ6C)+13=7bJA<2f]K91\><#_)S70aJM#+
// [I+=<9FIYEcOeF^Cb01^>.3PW9SGS_9+O6(#c/Q/B<9=BSbb?R@QaF,[WDY<ZeFX
// Q,V?LX<3(]@\c15FGM:b)GDX9+=.HZ(P37c[\LTDAZ5[J3PbH4g4+N/Sd-W<RYCa
// X@aRI3e<9/VJJgbfQLEYVGI6,5[e7<XA:91172W6:[VQAc>5.N[=J1EAIec3:.CX
// 5QK)GJ/9\K.EB9PU??W@AUQTDEJK?62)DGV^70B,_<EF:((P\4.CG-?H[[bD(:]D
// c#fd34Z68VCWW=OFFP53VgF3.TOY&:LE[HF]X=93d\4Z-DZ=K[HFc.Lb;@K@2;]0
// L=ER\5]JF]b.eKgb_K63,-NYaYYM3;7(=IARf@9[.2DOFR,4)/Sadc#K=(b[_?Z,
// g=D8NXP/R&9VJ4;D2:M7GC\W1D:e4e/DdN4Te+,3=BU=.8W8EIeL\28Q.6+PAY-#
// 7eX@[4FUDdKH+7\_,GH<b/^CM62;(VL4LcJYI5Pd>9dUVCeT)Y:P55-CM7/BT\d3
// 1/;/=D/4MM.c]9cRPU70K-.?@&8_fA=IdFdWBL^\4F.R(c5R;:IUI4Q+](fAKde@
// CAL/]HTcA(Mdc(,D5EQV?/9/V4.]Y?b?b6/E3ZAGL(U>P@B=WMI0L3?7X4LEO<9d
// ODVd(G9?UUg:;f&M-0Ye@dbfP<NQQ@&bfQ+e?J@C^X;BOWaS3Sg,fDC^U;.=gK#&
// eM);H@+T(]PM+D18AS3Z&RLOb^Y8_B1V+6=>2>K\]CG5e>PK:e96VLP4D;W+;NS5
// @V25D2cBcPg94b.-&^=)>HRS[B->?).G[#;#IWEY&fHJ\M]?K8MZJ.eSVWK>1;eL
// C9O&B0QODWFId_LSJHH4cFcF+TI:Y/]FMXY2\(^1(51=>-.c&C=D8a+6=d6&f]0Z
// 1GYV:<,.)3]OD8f0N@L,?gU1388g2>7=8FZ7TXSP[UM-(F4fd[6L4R56<dHGf=I&
// #1NPg\\+,W/UU+>JQR)bEC=,F-S/W:,[9D81H#>E8XX,B2U5b9F-)^D\^(c+^W0K
// E]+#7W?2TX)5S]:gFM7g8XS-&@_-K]D-L&C@5FU[\HD67Z#[L=[OK072Q@9.2GC8
// ^E_LR-YQ(9Z2]8gPfFF<^I@8dSH,0L;_CHL\>PSHW4<I#e+04P]\,Fa2G9O/S-P6
// 5FN_>ZRE=#JRPX5[=gUeJXBNW&Eac,(EG88O)I<Z6e#>X_QE9VA4Rg>QJ0aL/aOL
// >H]@8e+)WeA\1_d?f+/:g)0R_RVeNdT;A,2<#:WDAQY/+dAg+(XgFFN51F93C57^
// #=F\@[B3>@5\<5VOLPJ3@/ZHIN,a)gQH3=ZgS+7E1E,[f1E/077=X^U#GR)F=6+M
// [O\[QFa1S0A4LTDSS2]Z2;KJ2.G?4CKI/17?;CbDL(7@_-ZOQc,=5dL8.KIFf;/@
// _B932+QOd@ag[KF<N3C::[V/Pf#M_#/+:N73A8,M1D03bBVG;Gf[dM@9XeDZg[3:
// 4>A/.SBfU6T,EC,.DRG<Yc58C0e@><>LeM>1M:WO,b[#06&#HZ8b3([<#^GUU-FX
// ae97X(4URZ9A;VA&Q(fa;Yf7C9L(;FWFUS&:93LSEacf>LafFbZ^9#dQ)2=[7?>N
// NQ9)#+Wc5Ud>PJ;Q1_#UI+EL,W,_3_21O_W)&Q3(deS:\DK.4U+;A?:NW\.g;4PZ
// Y.CT0YeJ>4X:cD6OYR&HC8,,eF\/1DV\Cg<2@?;fTD^^b&7]fA&_F;TQe-fC]b-g
// ^\^Ic-^.MP(D9b<47?e?@_1#_b4e.gIZZ\-fQY2,:JW?KD1(#-HR54Y,HWd^aY48
// QW4\O@=+A7:Te,V1-CQ\0P(e-&T5\YX+/[Q,0cK8\^a<C9+#/EC_K>5V=fKL\acI
// +0+eG2Y=-\?YYU(?M_#/L6Z1Qg_E5gW[BI:;Y;D,XSPW4N&8P1KW8/fEX\,RX;ZM
// G6ea/QTO5<U2\5C4=fNY?C.-(7gSXGc_(Fe4372,23:_ZbZc-3ed[V\R+WgWEKd&
// RTP>E4X:MNd\83UY:)a76MQ>;d-WD:[B#F#+IQR3/KC.-Qe?NG08,H;c^Z)e[<E1
// 0-B0]c)>C4[1<\-QbVM/J<@XGO_d2=LRMcK3c6)UH+62)cOBYU[GeOV&R#+K#X9@
// dF&G,BZ3dIAE;K]7FJ/a77DYN3<^Q@&AS=EQ>K?(Q;;UF:3,NLJC90OeIR4#+VHT
// _\O/&?1X5,1&2H5HES&&;\]9I.,<EDggTB3e^2:CL^M)KD+bWYYcYLT>_US);&9:
// g98-C@0YL)?J<H[ER21BBCET2>TT#):55?0>_M)X,FD-gA,]S[,=a^KH44]I7(Q)
// ZY[bC7)N7LB&b+aJL<VC\VOR+A:T=^+;O<a>XA@HD8N3_,SNc9a0dKWX/M].;8&9
// a_2ee]YK<)dF@6L,P=ZJg;DcfbX,Y7U[;,=PY]6V7<<7<^K[=0ff+7<3B79Ff\08
// @?6RPC(M<3C9HR1G?ea9T1]4ec#9OY,DJKDSPKI<-Ke2B#?b(K_4NeSXKK<:dU1.
// :G=1.ARK\^,5)>S3/D5f)]_5b4D4AcV7b6J1+ENI[\[0#?-Z:/[CeB<:YDfS8/F7
// cc/21b_+M5AR_OD--7\4^]O23D>Q7[HTEOO22C3L19;VG@[<1BO66&6?WZ]?LHP[
// 7X=Q(@]5=F:R+^>^W90S3[<cd9#V+PG.=];?JMe#IR6J_V&a2)ag?8b+MMBe@_)/
// 4c:#.Z;ELEb/M2<#0JJ<cb+XRDSP,F(b#8_@FK(F37PD5K&K5:54#7Y(C[FEeb@c
// <WG@[a4I<3U[O5\B5R2Agb)M,FYaWPJ2PL\10634gQPUP8/J7<N>R&1<@YRKPVQA
// F?;36g>K#bWQ:S4[;P[SRfPQgeX23Y]<E>&P^H)LM;XDSM_-WGC9S/?(HY;H#Mdg
// WXXK_BD#Sa:gd[A73R68CJ2dc[V5,4BVGP++aSPB66@4C(@&[Wb2b,aUa441U1SP
// @]7QZ@YaJ770C&#6RKW#ML/@-<LP?80GT[MIeAG4OD)O6VQ8=aEcbMXcWd)C@XfK
// +8_UB0J)9BB=d-:&5b^VQ&Df+,(H_?f=#V.L4J_0a>Y,^9UKQK2,cH(I)]LAb2?F
// LN4#5RT)E,ES/R,eRT@#79H&N,dAaY4-M_:,-Df.cA\#H:>&f;G)G[+#M.][@fWP
// 3I\JSI-4]P,7e^+VD05+)XgEdM9/cfE/+EIZ7&QL?/]OfO_Y.QU+JNY#.IB,X^G:
// 830N_Df(,[=K]30,:C:&)?^CadD\)gA<H;EUd7Z2eKRgIC1A<SJZ^1GIab^0O/@+
// 8HM\:]\Q&GLTF>]a9DEWFR[>,G(,G@bbYb:[UK2UE0_+--<]P3=3eS9bCB>2&aEF
// 9Zgb4AM@;=K\+=I1P[<A=30L[9WNQQRJ4JRY,;TcY]]:N6)SUaN)2)RI:28b7/63
// HYXBb<3dKHEQV_7<aUM6NW>?UZ\>#_10-L><-3YH0\24+7B]/2dbQB.c6a,1]XTI
// )d,7a).P=RC0NS?7bBEBYN@B96S27YdQa0fMf[Dg]>W:59Bd0<GJ4SHWS4L4TP3K
// +QPd^^[D(=B<J99[Yc8X.JQAEHZ_3R@AH/<O5XPb=+b1@[G=CZHM3X-@^fd-e.C?
// _-eLDMd+K&OcNF=PePC^LN26<f7JZ.A68;&U,G:\2OD/TMf+Z5_^HPVRJ7Og1&3c
// C<Z?EWcQ5C-HR@-;73da,eK87g9MW:gM;DN]<<_c\M\LAg#FZJ/4fSdS#b^Hd9YO
// /O+7IVY=1/J:][812CD&4D<XM_R;Jf@#)DS2YTR>?GRfCQB:R,)f0Z+1\PFGVFIZ
// ]/e2GS_B,0>7Ad+<JVKbe+#f:==[=J,_^J=NE>&c;bBW87LA\]21AET8G-g)_/96
// 7eZ-eB&cT6Kb_VV)_7B2Q<_1VE(aHG6ebZ.KI<X-I\MT6\[J5F;4;^([4[47bBEY
// QdgH\(gc.c&.cRK:^AJ^54b.#34@e.a&ZW(>Jf3,cBAe^EdW[&[7Q-[gaH6OWK+@
// R\8G8RK1ONHa9c9C<7e]Q4bKE,cT6N_TSaRPO>_g9d5H:^R1R]KDMFK/d9IA+?CR
// AE:CCVG]ATT:U9e06SV.Gb7WVO[Fc@,+F&)(fE-0D\OF<E3:dFa0gQ9Ifd,bJT#6
// ?1Zb:aW=f)M.cTI^.=(JW]+FR2?HYbWQ\aBUZXB+Q#N>RT0P.cW@YSQ@>4gQ+f?3
// :WFBC?Y8gR8+42(2C:66?gK(G+;ES#O1>TBM(MeC>4g^6J1F/AT?64R9eM5PNJIV
// Ma9DVQ(]L_2/USLBAGc7>UE9\->8RBP254F1NO@/;4>cN4-6L5#KERPgZG\3EJU4
// JS_>A/77C+c02K7T=@+Kg(VG-cJTO#1RQB0#F,f=W_WR7#J.F>da8+,>A^RY3Z:T
// )a3OTH:94@42]L_LM\/Z\V7,]/N1)Q^:Je7J:/,)Z90<d#S:S8QDV9<57=#>BTEK
// D-Ze:Y@5S.U87P28dU>f^QTH7ZCPLH4W>BH^/QY#KXN)TQ2aXfPZRT\,WW1)+LM#
// &AON,<@HB-&GW]bPfGD_>OU3UZ.DUTSbZ<_TcUX\dG#b>Q;O-a\N6NKb+OWIcYd^
// a@,b5B1[SQ9d2I,TY2:<7Sg:NFCfCQQBA^\bN4EAF/RT)[4X>,I(<]#(aBA3&B:0
// S8O1SH3KfWR.SKG#PGZTLK^M\;QX&(<8_,c2?)>-/Y9[e_SeP5GAbY^Z/KKHOW2g
// +0Sg],Ba@_D:X/-NZK3_TE^XI+\6RGQ/KGF)eLC^3?76V,J?6O/@<T2<2GM@#393
// cY-Ac,9fE:a#BS=-X9cJ@/O/#c)&IEK\@[f]T9]eSU-9AMK_T58X;gcFV#?=4(e_
// e\90WY3A-_CG0+X3/Q5H>91.X:+2X5ce2Gb9HbafDN]VB>GP/-E>OOL@e6JaU#DC
// 9#[>(d20b>\cdE4#8,9HQNWC:^0DaaA.5:>MD3B/dRe@EK(#.cYNU(4fe2[U-JH<
// \>W/dU0?0@@HKSI1>6UA?7LaNf_J5UW2>I^WS(6>6_UbR5PD1BcYfO3Mg67AS>PJ
// CJ9B]eX=<TGXV=<NBZTL-+J;NU78]>-]D.Pc7U;N8T8M/AA>;<YG?Zf[.,0-(^,d
// g2gK(P=I9_Pd[[8M,&OQ@\2YKHf^4V;4/-/OD9G96M6.ePg<57UH>TC+&+_4LfXO
// @F)L^KKWCA6C.3fAA-XU08KUY?a-D/ZAA@-&XZ/d=49763R-,:NDO[cTN6dM0,S8
// >P0cLK2FNFT>(KAbb7#(cTP87U[SS[L5=N/\da5VIT#2\&a,,)SL1O,Oe:;ZU-TO
// )N8Z?]6CG>.XdO._HFRV-E4>\?BNTgMQ+&QCBM;2TQ]@Z<-[EHRgSdM5ET)eRQ+C
// g)Y.WWA&\PP6GS>&a80;S;M;]a..8R-eScGK@&aZ8)0LBJ&:^3O2XBLLHB9afORK
// .=4K/5SW6)#SSJ_(23:.Jcd9LadY:dKg9_;T6We++^0Q]d&8?G@LEOX5N9-6LcGg
// 4GfT6ZbD?7E^^c/2_=2eH):9?T90Q2-A#U0.^K_])K>G\IN>=UAdN^4:=I2EcD2=
// B5SaZ<P=g]2/_QX&>bUc_:+;88KC,=2-#AKM&(gZ0HZ5fYf:.>QY40^L\1[\MO0c
// S@7VMfHSMb@<R4,O5F;5)=B8_C&A)Q.5UGT7LEEWU1G8AP05M7\X_[R,WM0b[#?@
// E8FeNE9_4NIgX]?36<e-VE>f+bS+RF>]H2R8PI>2?0c,F^^C^>_3PT#f3.CR_S(6
// @@)3adK;3EG4GD/I>(._3QB-2K79@OIc8[W7,A/ZO@TG2-eCR5M?Fd23O_;>4a9f
// aE,=G1B.0NdA5>#6[GQXcXNX?BC-Q<F,aH?OcM?@<A<89O)6-_A?S&);0_ORW;d)
// 1W#.db8g5#-EY2.P25.cT[9<e.g[72VNDD/D7P(<fFE=))J;/Sd/R=ISG\:CaQ-B
// 8_\d3e\-@\/BKM^a:g2WHY2#@G[S&@4dE,EZJN@_HRZ?7>E:5T&;R1e?d[+FaS16
// EZP(B5LR@ebCU[[OQ^)f0VHE=@Q[(?^^&Y8&R>_=4g)UfLON/\;D[IU>TH85QBaD
// b5RPVB/2G;EeF_#eZ9H<^YKXD3@(5P]a4:W7d0;P9cCNWCKK=9F#_/N&R1H]TZ\Z
// ?11dc+1P(;d(TB-D8JdX-K7=FR@#WTCIY@Pg>/>CC,WKN&8QVPbaOf@5/f99GTAa
// 7;@BU8T=,^J:0V\PL[;^eT\;Bc^UCH&X]:b4;()2^6(?]THA\B9&+&/)_RaG5^;G
// OWWcKe[?-+gO9DDR:aMFdM,._KR51)_YM)UN8XC-)MIgTTQN\Wb(<B4JR0g)YV1>
// @2/P52:A8fBJF.LNE.R-E&I-).FWVINHWLO<K8EG>#JLF?gV/#BR;G7;QCFALK.3
// #B\6B/?1?b#-9/b<.?PA<B4>a#9V?NaL^;2T#bN00fGe7d6>_<.bAb;/S.K6GDe.
// QAd:FdN\(BTbTS<#:g/d;ebf3]#.?<BUfC@<XBE]]W5K3ZfO8HG0d]#+NTD<]+@L
// EE:[;V@]#G,GZZ2<E#.YP#_dKWEB&^S7BaQ:ALHP;6(J]-&cX<HX@5DebO6VY;dP
// d.6^Ka09>J;U71I)5]RZTeQPcJgY#6A5D_ZHa)-R[].;aE\a@UR;;8S-UY55#<\]
// <D&??2G)/49ZUJ?]24O5YD(5@?3?P]2P\P>./U1WMT1bK@KbXEX[Y.bA2=/\dGPL
// F?=A]E0:\\&\XQ2cW+d(+ZS>L3LT[HW4)RY7B(2TJ3K9eUW,6M,A5fC(HT4d]+B>
// LTQf@:LcKYY.Ec:7R.f(O/AK[0\gDH\gcd^>#M\05#g_N3B\]FG\-A)=^;.<B[NX
// /f)HKPgae9M^;fF-7bNY=&V5X6Z^FX7Bb&AY8SPb>CE03f#]A3J\K/.+M7f:T9=(
// UDHPE:)7>3@_W]\RV^75\Z+dLYBDA,.J8#,K_:D52;F7BcgA,#TBX0[:gaf=R^g_
// MT<cb7CDQ,BK^YVV00-2NYT5O>.64GSX+N9-ZLHX;?3<]MMF87eDDUJ^Ld#.<9>T
// 4LF_\f>S/SMK26J@AUYF&Sd(MVM\\&P2AD3_J#JeATWSZAAFXDMX>XWC<YTLX)PS
// LD;9:^@MN/U4LSg\\94.+84/58-ECaU94_B_269OT#IU&UcB(,g?8YOG&7DJQ13N
// F?B#ZbLWWNZgWR8QR+fGY0AKFZB.Wd41C.96]26A\X@\O#T#(M/42aOW_K3B=.YV
// <6BUgBJ:&T]DD]e;F^(KA(CdAYKR<.E,0J4Qf]R//F4K1:7&V,PB8X134FY?7#R_
// _.KVZR9I00YgXECQ\GHZ/PM_aIEfN]=@-GOQ92I[ZeCJ4T+a-Q-?WO>?-7Y;,XG?
// .EKecCdXYWLeOK_4_(@.4TKDYD(M[=M;=(XTI[V&7XS.?^GfS,T[D/03Lf3IIcBA
// ,PU^b3^fJEO@@S.NX;3AKCUJXZ+_])-J.LN0+.)[/\dN<dPfFa;K:ZR3?O.d-F@L
// -0A9@L6==C(2LJ1E@>Od3+M^\0UY6&YcC=\H;cB>8<5,+(P0=7A:<c6Tf8[6Md]Z
// MVA4A.dZ+f_>K_C9G2^#2[@X]X,C29JGH+CUR-E@fMV6HXOKKKH&Y0VS/6TABCKc
// (T6=K>d2\)4.c,:YXHI]9TgYCO\7CC\LI7A&,LcH\K6U\I]cV7=D/LX-\O;:Va9<
// T<GLaYe;&&6HM[2-7N;IX4[8g3Y;5<caQ+BaK/\WMDU:Z_fX9[6Ld7[-8d]?b^.d
// RVDIVF:AW<+7,<X]^f5L^F2WT1g<J?4BC>gH_N#]@(X51C+,ITVG-c#S<9BZ>dK8
// LY+-0Wb@aeOM@.A[bCZL9WL\c2PRF)]]7@cg\)K<P<[W&=b4]<fU3_^8ER6B(L[U
// M1J^4>H5Mc>&2:3JQIS53:>6R867W)bN3A6(;2H@dE+a[=M.fERH?8X=Q?b,2P5c
// &^>6#HPNBE<XN?(#gF<_WF2)IJV\I8/L&d>2a_7Y3X2ZEC._SYZNE)O&bU[,I+Oc
// GZ)])2dZ2#1&eLD[3(MHDL31SYJ/[8QaNc#Dc?;6B(3DDYVW#d5]HM1?4.1dW4SY
// #f62+LJ:AK_18Y.M,5aNZS@V9<Afc,BNLQVX[T1e1aF/09<JWEd&R/_-R9ba\JZL
// eHK-5bJ11/WM)c5[5Z;2[V0E@02-+ES,1#,,]4Xb[aXB5;Y77+?/Oc>K8HAe(3Y=
// TO^7IH5+NHb=9f?MTaMFbHQc+_S#=\Q[/S6b37?9a/:4SeQ7)E?25^eRLPPg5a+E
// 49JQ8UW93\@IdI@TU/Dc<;8X)/:9,(7g#,\/8IfP(?eUEb:7-?^)6[gd#Y&EHZA\
// E.1QCOQK]19>#VK@6C@FfER4Sa>RffN1WQDD6g@>GTL7R-#A[AE/b^;KR?G#F\CQ
// NZVH_Ac&ZS+d^4&=-Y<46c2>#ODS>S;4_f\EcaVE:+dJ:gcZ8-VfPDPVY1L/#dWg
// -(ZYL0-]<RJZFdM?;;8b4(R0DOgV4?<6Ld78&;I.:P4+LFFJ\X<#FS@f[]0E8b)@
// -45]6>E.@.9:59_<ZM#B#bHeC>J=<O:/2Q,0Q\Rf95_:^TW:I-Y9/?0XSWD:-11U
// ^#AU=VQU6WE>?Lb2LB7&F+I\dM1CDc:O8b+NDS^<#E\H#f#(DM8QfZ<FK/HdOMD;
// ,d,/H3A1W/J<Z&3(d](\Rdf&@/R+?d;LPK>3QA>U05N0QDab.GBDb_I[@V7CG5Z?
// CR?>LLMH3@gOKFIZTU+;9RaK4c7(G(B](JbJFVN>g9XR57TE,#227AcR^@IP>W9_
// 4gWEKSUIUCcRYRQcB]2BWZ5]QM2d=80=+^IOR7aG6)@7DHTd0CBVQB3Q6.3Y=G2]
// =6V^R:JbXUPP)LHF:@YZ)7#gZ5cHR6P3=H_M0^MB[VgB5T/>\#Bg^IJ\./;@OQ.N
// IWTO=?3aPM0-Qb9K&-T4Z=0Z\/PdX?K=AY9e3B/#/VOaHaIF/JeM.cWT9\2SVE2f
// ;8RPc2+R#K\Z@W5JFFGAbA@3-aF98@9?D+705?T3bY@2VE5c-aRGL/?55IJ05SdH
// BaC98+.IU6>#LaJ@ST7LVXS(Ag5WC7@&ADaF[RZbFD/6Mb=MWU0=WO?<O_[JT+/&
// UK;H6KPb),Qff4K92HHF&bQ1&0.&ZcRAB@]E@1F_^W<(]8GN=C^Wa7L5@bJ]@7:(
// UA(;2&Df4Sa]6&^M?&?V+X)b-6)T>NBgLJeaDD;YX-3C/NFa]^5:MLAXc?G/0/fO
// a_3\@UOWLYJd-WAE0bH,.BB]eO@^WRNHWa_-.)2MKW#gHf@\\c10bB7fS:E5B7Q1
// ^?5WZE/DZW4G)HL;,2]MR>,J7;U5S&:+g]Y1,68S#B[?P43-/?^R3/FP(HgQM)bE
// 0e1H./9H4<M.AGF-J;B,AHW.AYJ>A5gNA00#P9ETQ2DPSE1G4_9][)E)5aa9Q#M&
// c:@YLJQ5RQ6Mcc:0QO#9@(3;\?\:83:-Mb@Z8WF5N3R)Ka&L:ZV,S(;M/d.Q]:YN
// \aMN@5>eFcYIF\(O8NNO0g#f(F>\D-(28Q:?I,ScXEEV_b0J++aQ)5<5#QA]K+\5
// )TW\[R.^NYD<F=73RdY)gUH[Z[0VEOccMXcKXBeHSB1?>U@C&5D6W#/OSM?NZ_fJ
// f+,[BNHX.Pbd;c<]3U)[9U]dNMO&Eb9GNG5):1O124(CTCce,&#]ZIS_]JdfAB^g
// DEN>I(,;[WHb[JMLFQA@?&fTdZZ_0;@e-94X;b]_?[[0A=I#)gA\O,JPMg2[Hg\B
// :eLC@B7,dDCA#^<5SE6Z+M)+UAJ5S;RY2E6Z\@]L4X?4:g1[#XIC#I./77UgI\@X
// [X^EKDCFCOS+Ea4::G^]T2A&F[J=I-d-G,^HZI:V-ga>V/<^,ZNX^)>0P,YO0Q1U
// D1>5-JPRVQK_EKbWXKB;?c</]>YPT4d[aG4PNI3beW^NZ^fINIF&=90P\0I&?N,.
// SN9Cb@1aa[[/7=,.^-_:+?T2]-5<b0N>SQ8Z1S:;O;[E+/H#1]+e;36D&6P&;OAP
// M#2gZ7c14&?N&PbF[b:?;&;2gB#ce9ON[LNQK;FXSXV0]<6J6MYP4U@fZJ9f?)&#
// UC?=OFe,N(LQP]U5>YEfXG4Gd\79&>6ZKZ4dg-@-B(:.4XE2KT,<I+6eb208Od\_
// [c,)#L8]a8B);fAP-3->+P3[Q=<GcNX/e+P-K63#>]be-LbXN,\6Ee>C45fY3)W?
// _;E.7<]N]a7EW@B[T2BaLRY,/cCaZ6(dYT8=:O/cF4/],L#e[?Ra0M+L4f<6Z2FN
// C?[Z4C#(Y)0J(+b/AW)dH\;/E636Ve=bRDO>>e/Z_8dg0/@_=G#gWea(>O5J]20+
// O1g\Bb5c^/AF/\@M,&88QI@aYE=(\FUaX<d3M=^^2;:6DG_&VPYA2;P?+cF[Sa>Y
// F9c@KW]QGH2^Da5^1QUdXF39+<a^JM-dbe_WQE.KddfCVRec9(B8.QAAKU]&9ZK=
// L8ST=UR+RJ.OdO?T6(Z1.M[Za4gd44[JQg1N@2?U>]G\)Fe6bWce3OAP&\+PUO^C
// 4OW2FY+:Y6S.DP#>T&S+W=7R2AQ-@<C)bd1TfI<TA8@c3QQL&A0\dG?3ODJf:e_9
// S+\bZbSf\.W^ITLUGZO<9W8I,4J\aN,.))>TXR>,R;)#T+(2)=S0f_Pc4YL),4dV
// )3WG&213DdeX3T8aG4dIP72Yf\(81M2@J]9[[6@:7LB5OTW4]J0>=,+DT/1e)SYM
// J(dIO;8LPf;>OY@Qf@?/Y=OWVf)cFZIaFDPYC2SL>--H?^M9060+HER>4VV?SSd=
// ,:RIWZ4KCB[OJ0_8:F8<A43N;Gg+Bcd3I&?T)]K0c8]S+:;]M?Z+5VRQGbJ9)Y-?
// SSeNVWeFeOF7PJC&&b5;)R,=O5[f34ZQWS63+d.ZcY^UK7AQ:>8,/\AMUU)(\-G2
// CgeS1@#dS2VdZdDbZ=4T6#HaO,T-bUS5/.S&G]@P04=)KQ6([W:=QKK+?W(:N=Da
// gE;fRC5c5D_6KC22fgf9WJ\CDT66OR+=I2YX2>)Z2<a,Dg,_9PT_FaFG\YUH+ec&
// c/df]\F)0FU\0U1aYIJcR6,>gQF\MD6#Z)_:U:BQB=a1YK?5?,,109Z01;V?;##L
// FWS&+3[6eNPbY(;87:0Rgd\dD@G1/FQJE1_1,7:@@UGe/<:^96-@GS/L4I;7Z3=X
// <RY]c9I_YMIFK&fDdSLV-S<gF.2P4:Z5@6SDYP4Y68gH]PdD@ZOG]D(,N5UCYP87
// 1..6_>)X[@4D?c4)1#-;ITG2_<b=NT#FWP<5OSS/S^EF)HC=C6SV(L5aba[Y(+D/
// >/:e(RNMIXN=HA-eFC^;JfeE5G6[LE;Taa?7WbT6X3UBJWUb]FbWTdY=B(J1R&H=
// 9Bg(7SI-H1_CVbB#:-I?g>NRS\S@C,]HWA>bSTTbZOU_;TZPC2>CP;+MM,EITc5:
// MeC=C596TaDg7:bT;,WXVUD^2A/KBUP)5b(+Z6;A#&@Q]DVOH+?3H0T<D;gPS<KT
// :J^S6?/]4RMD-9N\]-b,LWQ0\gCX^DFV91.@>g6;HR=#-1=cPEOM:_TaSJ=N\04W
// \^?^Dgb0ICHf5a)CcWBJ/Ha>,-2N^>C7+=>fA#Jb/TUV;1CSdNe0>^QP([0MF<G&
// d7)<RQI1FR#Q(-aH,[9FIY?8131=/TSN\E>GQN@2MdP#d-Z9&14+>KKB]]8DK^2S
// 6daaA@O-;K;S8GBZ[N2ZYJ\=^3fBZe+B^K^>__]9QgeQJ)WRO&1#.^-558TCYWf0
// 4O=PG-f&IXe-c1Qd4=aV[\@NDX.4[g,CI:O<dK@@)Lg1ZW4/CCacOTcXRT^UZWZe
// QWa8.c6R[./B:6)+g:WA9TYC75]8F39>^MM)G6dB_QVK)WR#<1<3&J^HSRBQ=[c)
// @__)(KXbX:.9+30Z,B16TN>IAZ,<>8a#6[#[G)Yd_3W3Be,](F(4(d4S8_83-7;e
// a3PNHMK7fQ.9MdFY36F6KFDE(+Ec>05.4A735aGbcHZ^.1T_NM\e@AN;Pf^DY1CN
// 4]cP-b2ae:TFW0C?VS-Y;LX-N;R8AAcH,MU>CHMLTA^,[D5KSNT539c-ZRUS.c6[
// ?1->+1Ub,7.Ha26GcPY)M[Ufc:5d6S<DRX:FU@XG[=K_5R7J5dKCYdeSK3eCLOW-
// 7_UO]5&^12M.D(<W?G@<^_R]D[\S9RUc+4I6-^>cNZUPAUN?)BA#P-?>R\>,de>S
// /ba4Ha,G[[:c.&SR@6R=#VW56A8gF3ZUg(,89e66TS.=Q6]a)_QfDF1B_XUHGY9@
// -RcC-)WO>Ce3MM)190/,6R2[1IK@JZG<37=7WUZI?)X.8dKbb4A9C,0@SPe^QC_=
// 9)KA=Ce(R8Ca4&)EE7eW5YGDcK_+;[HX9g;dIQX>fN;Z9]>Q8:fJ8M.Z_]QLO3<<
// b/>>0adfTfX.YdH?/aa7Hb.f+UPc]P&&7\,\G<F>S8;Q,YJ6G@P[\9,CBORXg\3;
// B&d(XU#:Y_agM.C2WG4?K6_]V\E::D34K0dg8Ecg9.X9^Ofa4T,e_BVQE12_\P,^
// :6J#gE>U-;-&14UNaSOBE8,^<+.[4QNIM+?QZ3U@JL46QPB5VX9J1?HS]_ZUM1d)
// SODX]EL\H2;@47TI3H6R6O:^WMeU[U7R6@\8WA<897;=fgG#Oddd_WZKN[B372cA
// [UI;COc\6;\2L9>_5GH>B7^b+<@,S^PHJ-@8+0K2BSdYZPO4dI4df9fCCZK5KW0Y
// 0@b+38#2g6Q5AcB9/2gMEA)=e8[GU9WGLP9ac<a/DA8N73:T9PF\C,KV)W0;M\1,
// \=Q+f]1afM>fdf];9RcEHOKVO-O=S_=0&,P.LHeR@ED0WFR.X3NGI1+NK@G[YV]@
// 8X@<)4HP=#//-A:<f_,8&c+L<O7M+5]YEVX5T20051G&P94DG=_,83S^ZINNDRcO
// 00HC>MQY,=-,gF:GTcSOXQ;Z//0V8C2>UR^26H12=09_OQ3N5NL(G42YM6)?F;.F
// &g5:fL#0Y<g;1;&W=TWU=J.N#1>F=YMHff+]C]7b]E>Y@ZPAO#ALL6+=]S^IC0#U
// ,O9I9:P5HG/X6M#0K,2R=60CM;cd;A8A<Y1?-?b_Y/XNAIgW_)6a45M_&P&),0+?
// 4Y(dB)Q/H:(_2O4Z&d(AP5Z.8VegE?NC_R7:d8[75YNFMSbA><Ud:S9S/8.@c2IT
// NTX.:J+;@ECKM7F\N^GG6YW5,;1:U/aAZM+SCILMC+HY,JCC4[e^cMA@2J#8JDcX
// 6Y(S0HTFF&<UPc&F9[NN#)XB;U+3L-CZIPZETQb>V;R;LbSfGDAaOJ7Td6/f\=:<
// ,#3B+2WO8&;:f^;4,M\LbW,NY^9TbJc>^7C5^2d5ce6M8IWgN^dNC0[<^4M7^]?(
// .C0FGT+7#>d3&3&1^fe,[..\eVa)&0.[A]a+;UFSD]d[>c]:K1Q3\XLY,S>b^W4a
// )Ja+?C+ST/FA)R[[K/0KO-CZR,&[SJ#>a6c2[TP]9<;TJc2K:]1RRFe:U?;NH#e5
// :3A4>SBaSW5e]_5[WCL/Gdf[PU8PCMLBeD#9@gG/bL0#USAI^1;>dW+J)KGd]B44
// g)HIM2A4L9=P1L3POX>FZ]CXW54OBb]Ja^H593d.Lf5J,K#KB8+PD\bK>U]BP.-&
// e\;Fc8B.WNI@g:U3^MWeE0GBRS<?B&CE[)5\8=8cd274&?ZLQ_G4\9CWK9NXQK15
// ?3FdB^OU5(,aN8-RI7>A6R[5KZ?e1Jg2@7Tg6_5\U]TJf:]FTFXEWdeETM3)^?17
// &BW5Z_=P.=XAP:0;[KaGCP4;1W::2\B^A\[Yd-8OP9eT7FJaRaH^gFJ&ZHbSU8aM
// \=&ZVG)Jc?SG2EB_(/OA-UA3]e<?63NfR/(N4>IKd#FL6#7;eB1U9OG:;a@,RE0T
// Q#UZ^NJI.4Z[Zff#S<+K[b.E5aR@AGTE6<61_0LbAXE6.-fXVPQKA)/bP@#:N[BG
// DXH4_;_?1]S^^H04[RWa=MOKT?Qd_(MXI<9H7[5(:<D()eN9(IIVEUaBV)C(-@+C
// #2GZ1g/O<GFPH(R)JPWa9BC0BENEQ948BdIE@6WFBV1P7GE/R6Z;RZJ+K.[8c#M]
// AO8e9b[>(N@:;:8Lb=#@1E:;cU\WZOGF7eLb-L1e;KgV5CC\AYZ6@<M0;W5N7;<K
// e==>3K.]-+U<+91#J\BfB/&<<374TVST/2^(>b]0OY^UM2LF8fQ_M_Dd@#XRKYB)
// :=fc]ZHK]13O-,N80_NG;He3e4VLR^,,#C,.5[&fJ\8K(3FN@[4-4P;NAY,H+^aF
// fbX_TF(V[D9/.4KTb4:+8W3P32_VYSaG\Y?KHQ;9[]E0#40GR.-^.MCPVfXa(:ZM
// 5FR_;J)]46cJ[d5>R^WY>N&NTNd95@acd=VE,@FQ;.+A@-GJe_A/<6bGD_12ULJ-
// MA90)>CA/4TegW-+0FD]]8I6=Hd^E3eC2g-&afM?MD?b[89<QR-WI?K.NP8)@(E&
// BK_=d+DcJ7>?-8eMa[N<QRMQP#d#0POFE]KK>T_J,?<(THZad,4gHLGH[?>G)0f+
// 6a^VgcA8cUE\L3M0Q8&.ODFQ-#W,JUMfd8fRAfU55W1ZJ.G3fg5Og=7.<4I[[QLf
// L4abEMHg@g(WP#W-=;e9eZ[<^3F\c^:M500O@/[CaABJ::RG\DWQA)\FNSA6Q1Ge
// gQPB<QJ^RbT[e@X,aN/D=R8B@JI-aafII1<[dEU04=Q:2=AVb2beB8K#N]JYM]AF
// [:GM7e?R:f._P21C&AO/F0BK(ZEecAeGTG283T<;US#]@<Ae9Z-1Q@06H5AdN<Tf
// ._cBY<JVO0SZ.XVPEEC6+bf&V5ED=N-?Sf^4\Ac/V>Kg>V6;@B(_>Ne@Gfe&?L4Y
// 4B>W7<TP01S_&3Y7.I&#D94-cUAF#Cf=;TY/6D-\bQ8dF2,8#4fdaI2@daXEQbDa
// X9I<]\bCaKH[XJ-7FBH@=)@Y5g<6IUXCPMW_&#]LFDe(:<d.;_Y1K9^K7a>?CMA]
// 3?MSdYMgbSS4^_3GU\4.^<L/#FG:;LF>8LNGVQa7:JSXJNJd)]S>I2/I<NLJ4RB/
// T0]P\9bS,5M;7KKaQD9O4ZF@1TD/f4\BH6<B[CU5?/C]52KeUOY[eH[-8)#Y;/N1
// MYfEXPgWK8cSUEa,CVcGG>0U7V2aX_Y=0&.#NZ697.Va-cFLW>4;S;>0X)Y=\:L7
// K/I<B2Le1OMGd,O3O2f9(STQB(,eU^@RYcD:9,GNdG9Q6>RcF+.\ZQ6P,G<0&+I.
// +bO0f]K;K.BO)O/d>4R:]Y2g4-FgY/?5b9PJc6#,X:.&f8HM8f5.QbR7+ILTZKcU
// 4G\;5CW76(+<&H-W+?#\PC#]Nf&WBT[:6IGc)S9)\0S7VM>@UWc&N]V&MI0_^BI?
// 7RcaK&70d:@67#NG;@Yg0;Td.4I64Q9G>bbPA^bB35(9;9AE+#0(BV=Bd73^GIV+
// QP1SV.UHD@dRR>U(UJIdURH]dP8NU/<U##H.8.dBb@SdK:[7Q=1:&]@4.Q)^;,7L
// ON_J7.TY<F&4BdGbd=dKe;>^_b@MSD07;9Y4XGXK386;gY2MCP&[L5EgYH[=5;dR
// \_SU:5c/3X[gZ.PB)f8H\0(X7DVfPW6<caQ(.;M1QW,@KX6,SBM707I,#C4>74_9
// Ab4bFN?]O\L[g7@Z<f194E6-<(HSb,cg4:-OGbM::\Fb(][_+M;Se,KE.I8N>BXR
// LK,A28g[aC+c(,a&\#M?1e.a139UV]d2:0Fd))4f[V+#>_W(:g/,Y:f[bK;Ff?XS
// T2;4:Jb_I8ITfbIc0@-eSfbYfQJQF=S=O9&T&eWBBD6A9+Lg[QVJbO^3b[6Ya?1)
// Dd,O61.3)4L5fRDb]C6?9/8Q@7.SV4W>4Vf2T^:H@U_e3BY-]d#Q(^#R^/.,aD#W
// V@aL?[>@IG;c;UP834K5\PfeB=NHSe4;EfN@OJNR?KgRIa_1F-H?80d\?I3c_P(E
// a&/,VAABH+#)WMOeG-]8@Ng:7ZO1gIJ&cfR>#B<W<T]UL[6ZY(Z3YUJad.d[d-2F
// a6@g7dIfR:OYT7<UZeJ:TSbH?#V/:6E?NdD(K9b8FHP)XXc4K)&gM)Mb,1ACW[43
// )#2>U0)K[5>:@8/.PM7cR.JIP#M\\(d6,-<bK<-2\8/Le;dAAG<SA@K,)Ca24EXQ
// cVXG3[2LbfR@N,ICc(R@N^.P:R3HGVg[1M.LZ/LGAd[RaIR1gTE76##BED>]U6X-
// GLT/cU]JRZ^57)cJ6LVT[4SbUD^URMd+QF-C>28[PHCLRHUA6:f9+a1-@a3CCEI3
// LBe>]&-)e.7?_(/dM8]]NEgP,OY4XQWR4Cc3T6XF-3Kf_]9B_:I1;e)KVgg/9SJ@
// JFNcCS7)K5Ic<M._@)8J\2OLY7Z]#74HWeH:GDP\c@@4(QPHY[>>7OL.;da_FU?^
// ]e[aUQ[d-MdU)\]P5\4\6O8gPZCd]>:&QBM50O;/e4]UEc\(L/N,@?B]:g;N)WH8
// 8D8(P4a<Q<A6EEg7A;4GW\W<\JQHcAQF+]LEJBH#7:S+L]e.La<VB@VOJTGbFbN(
// -ObT9RY:ge@FaCN(Yb1g5#_^G,O\_^UT#fa,\=2(2:&/^UJC]X]3PE.Z)3Z=)#F@
// g-T0_#YTc6<N>&&b@c8bX^0Sg99Y:B<BWP#5^+^O#2D2_NU]01g_X)Y:<EV9S?4C
// +ZFFX[/F648O5]HI#NBTF]cXc?^efRPBX_c/0]&/W?#,b]-2_RIbDC[HW@[gUYX,
// FXN]ISYM/)e.<ND,F=QNFM]VRCHH-LKSZVEbUG]>Ib8Sc6,LP2YdR)[d5J4DVg3O
// KIbaY5=N_52:XGe_X-I=)\,;\J+_c>_<W+f^E@XAS6g47#9b)0D3U0G&8C7@+<gI
// AI79T,^=HE6/TQcUc]C,Xf>GSJcGgeYa6cI;3+[F/FFDF;Lb8V46XFRW\?]0c?1;
// )^EA&d==^V9_E&]N#4I<<E9L:^?K]LW_)BFE@]7I<EJJ_(P3L37VfRaJ])T0^IKS
// =\EPb<61.f/\?LI524>?UI?5eH=IKW2S\;Z#,f14/,3IK]O)DZ.=D><9LA2^K81>
// >YMAP1@\SMLdIHLQYR=<6gZ\c+(eLEcfLC2?&Nb9eCX-PMebcTONICC7d1<>@E4G
// [7#XXB-0TNT^)Qa+_[__&8&5:d7.&:aebaPV8I\ePRD.N^c&JBR2S_4O5<N-&NQ\
// U6/b5#&5bTEbO;54Lf@L#CbUV/4HI;S<D5>bX77da][LBf)<N4+BT(AN^6NDGg]R
// ?GI/+IV#IYLZ^#I)YYXgMH_GYf@7FDNWP,HT)#SDW)6Fg/-+O\5W,S2?]PGOIU8R
// &HcNV:A=eNT&QbKc=6#_;6PA?H5P(<L=KJW(V?&R4e)bU?V?Wb?::UB2MW/bC-/P
// X3d0?Z5P=/#afffdDB-00babTVP>XcCT?a<PWRI/#FW<)3-SZS2VF<<0Dg;ZS8XV
// VKf7[Q?WEAQ_JM[C)G:,@;R=YUAHNK5<)Z.G(I?Tf2d[aH^-&.0.Sa>7D4C1<1X[
// dRYdg:9L7(FG]GMQcXV?;USFP^&TJc7f]B5KY+Qa4\NA1\GM/3T/H<1X-60<NgN-
// a]?8G9c#ObfL]RU[E:fb7/PZ<)B8Q+B&>(<^ZBHa9W::N>fSJ.Q47Y3&O&Le:0(O
// U/<]YH\2Ha4RW]55XXB2[K<^.e.=(:@->NYF.O&&)RNYfX[75._0&)e02JVSBcHB
// J,Y8S6@6^IVL^;&Yee56_157FQ8@fC..+bA+V8-L>\cIePdP+T6@B]9#&]AIHXdH
// 79bTWZQ+1SbL&CEG_F)-+?&J@d3F6T3753=aZ^aQ.\L[ZZGE^7#W8d=4E_TQ86W^
// 1L8Te-A3NU4^b7)99e.H8=1OV@K3DJV,dZZ@LM/UegS;8>gW^[H^0g7#-8M\eUA(
// 2EZ2Q-:=[Q[W?YE/)/.J-6MAREB<f^FB_\1LeI?IdPTHDIG]HM2H[#Y:F5\eD?aY
// +UL,TW3-E3ZGe^^Ef)5J/=GLGcPT6[LI02TKTQSGF8a5@SO[_@\GT?eXbg<b2O(X
// bB3T+O]FJCg^K?W5\[:O>LX;8\<bP&aVBdC8aZ;Xg8B-:e4L/FILB[@=4=R+CLE[
// gH4XDW6;7P;VI0L_RGa?PcQb&B,GG/SE9+Yd2C+0Nb-4e0bfZO9gEQ>4>UC9CA;e
// C[)[29U2GU+DdIS))GaRD\OZMaVIE(BQ;[;=;\Q>BUFeA6gW4[3<JDI/J3_a56R^
// 6<(eVREJZ9?]F,;F0&b.CJXX\IQ>VaGR/1X>e#1dRQNfeNN:Q#?F?3=GNFFPg:Va
// 7+FJ@5-L=[]I?]ZeY=LF05Lb:dOT45(3\C+gKCU.AFe4gXE-7LM85STe#J4UbOW=
// F5?4#[AgP[#E<)^84H(2DJO85)f9]f&/OZ\(G),+<4W55^J3cHS02a6+DFSaHQ)6
// ,cIQcDPQ^]O2Yd6ZI7:_L/9#c+C<NGDCecDF@cCKE@5/MBST#=-#eRd<?2OPcVUO
// 2K+@GMIN;&e8<M&BAg:1DZ]I98BP?-.&]aTWb9d<:33f2GRL-68Q(<e885\N]9&]
// SbN7e[^;:6E<0(dE9P5MSWfOa+S5DaV)Ec945bK<:]#07eM5#eOd0U7G(HTAb>Nc
// M,>5,Xc/d695L6#&.=+TNRZ]b5PW,gV99&AAOAIF1e0d&7W7DHS:^CH369)26J7]
// /a5Yc47eM20;aa\@WL?Z#?<OQ>e-JX4dEZ->C<3AGVH4cU1GCYD-)Z?+FE6&5#\D
// VG-RQ3a-W;(?XK;G[]PA7Ufd\NP(<SR<)1D5@E79gg)A]db6P3[4af1Q<A5_K=#&
// D+<6HWEIYZ1E)&D3_+1A/BT7PJMfB9DN.Z9;OdLec3[G\&-5;ZIP20ND^>cL=Tb:
// HUcKMYS41G_IcA^R\PW^)=dPF.J3_DSSJQ/^^#C][&+K&U)@^gU\@7><De3/GF3>
// WLO9+#DVeQ<4g2TNOB6DgbG3dJ,c4;M26DI]F:13JNZJe3,bDT-_RW@/8G\)G@0I
// ]AX8JM1(d6W>6D)MYQP.TP9GT#TG1eF7O9:c?9RB[)B+<V14])F+G>]=]^(T[#.-
// 95X]E.UbLZd\ZZK5KGY.\^e?_?R-Sa#e#,G_5@FQZ#cfY&J<gKf4EJ9X/dY^2eWa
// W^(V<@7W#T<ffg58)N)=5W;eQ@:=J8RKQ-ca)>..H)+9TJ3]EP>AKE/9SAY0TSDb
// 8WZX8&F-_ZCM>HRK.O#V:WQ7U<cEW5GE1U-dV?BO]bD&E5YHdWV^@35/Q@4aQIJZ
// f_Y_e:I],B1#J/aI&R>(CUTD0?H/:ga^gZRb7)6>JAVMN4XYM0a&D\TVWO,3\^Kc
// /D>CBZfZCYGUM]XQ\Y>BU^Of(Y4#?=L?.HD,_[3,F)[]8=K#YgXfL]53GR=De]cc
// 1\FLSXa6CNM)AT;dW6B@6c\#GaEH<#-6)]^MNA3DX8I+cc(6-fTBe-L<8&eJ:;3L
// &f=Y3AI>F1URMPA5DNCZ1d@R8SR+HO[0d3#\?cKSEO6bH@.F=I+,&UWATZ;c7_,]
// KES7V?)1M8N#M07)5QRSK_=DS+7G96C2JY:FN]&G2RZ]QP8LbQF>B(3^)<O@3<NL
// 3Id.D4TN\[TO7?C-e(NCGaKP)-3KVa3WdcbX6@PPg(MI;7JKX400aB.?3D6CfCf3
// VATAEX<LaXEKAaIV9PR]UWAYa>3MH?eZCXI>N6Ne]DQZ,R<UI=\F<_:25A8aCE0E
// ddYWVQ5+W7W-[G?P;_X.X2(>#BK<8/b:T-VFT2]J81\b)B<.9g8G9M8YYM?b@S.L
// Fd^?2PUGLFWUP_2>Y1YbFg8:/f6WgdZdd@)34KH4SYCc95D\Qf-[TAfBbPT8P5^K
// JE<P:bM3APc+4MO5H)34F;JPeV[+dS7<HYE:4>2gULJWd<F.@>FRI09d@08/NbfK
// _YZb^YL2OS=d^S4T9UELMC7Q&&.KYE^:ZD[YU=WOIHd,[Od(9L5?K0KGF(,A8BP,
// 5#+^DO.)FTGHb3GCFg4g<d@N\c2cF3g/Z0QUb]AZ3Z[_f;W2;7>]32\\:(KI2VN.
// 2gF0VRS73@PF^1V8U.^8AA>]gg3^UGgP#I5:5aU57^EJW\L;TR.JE/>FZRM)\(NR
// AN++J^60FPRNgFC(#;>Bd5LNIWTT_FYBB;g85/Y<U=NYD(8M]UXe6.N6:([?/^-K
// eeZ(#-F#b&:D:1#)#F/FT:cP4F@Xd00cK+a8=;<QT-Xb?GA0&M;Ibf?Ed(gKU7I#
// R3\RLTCADH&AU4b1;d8fZUG.Rg+AWO5\fJK6QKX;adcN33VP4e:2c-:MR7=gcL9=
// [D<9cU<J9K76BU@##GJ;g5K/@T)M]AEOJ\bU3gV@NB@:-+8D&HeXS,X/f]\5-IaN
// 8<];[#9K]\(E_:EJ70&V[TP5^Z+QE)23P[72+C,8R7Xe9))N?c<g-a6W^-HTFeV_
// I9[+-ge^,2R;f#71?B)[I].G_CXG\)T=EUL9>1.-SQ5W5KU)?B?2MfY0Z)W2DUa9
// cLccbaf,QEJg/Kc1\2S&L?\e:-BcbHP#@<(cQ/0-?8+-fP.)gZeTWH_4g\HV79f^
// (c6?U9QRLJV9_@S7X.:2^g0=R@R_SBOOL^>YD8aWc1JNVMNC+d?]ZT\bG?FYE68D
// 2+7EB9<ZL^-=B7?EX;dI\[?U<&=4_+F=4:OeLOe/=BK:Cd7-M@=d@L>_/9:AF&K,
// [3;_B90<WCHN6^O4#[6=2.V0VLb9^ISfG[_>@A(EN72H#dT[]e_5Ce)8Jc9V,/-J
// /EaSK#R-=)aP+X(L+dL/J&&CfPQYY,E@?(MXMA<c-+\G^ZN]6T0f=B;K43.\ME12
// #H)GcP8UZ4gDa[]9PeSA^^;NQ369-MP@\UX(,4A#97@eH0VZ/FZ#cH(6F=.C:-8W
// ]PUeIR]Db?<HIK::2cKGU]?/]GT2VR^Sf&<0?#VA?.F@Y/c=;NYA_J.\f>W^+I<E
// =d@IZU&@WdA/\e9)Z3_]4,Id[;YXL9;-bXWCACCAZNR50[QM9He41,deR@3V2X?)
// g2)S,>+dX[T-PISGS@Nge2>+=^&9&e0V+KVb3&L22I\9@U9-K<\I^L3B;_/X9J9T
// dD7+^97CBS2A;eK3UI8d+SJ?>KDCXC_Cd6/d_GK1LW#R:H#?G_<1fA/&PXF_<M[b
// 5ef@CD&)LHMEg+c[OR&Y)0:b])UI6\cL(9gPGc&.A3/#A;AHcVKN.C1T_#I?d.:V
// (]@H/AS1ZDNbeC@7R).N/?e(HIFPW?8d=?H)U:)ff=MUO-a+BMDA44G@8FIQH4\d
// 2-d.]]^9>U4>72OQ&+?DTb5HYVQW=-^JQ@a4FB;7/+2>(@Ne=</9He,.CK4+d-_R
// TC[00<Z(MH_HZ,_U3_)LZ+#L<aZ>Z)F]EU8cN;V\GdY)Ya))SM4LAIL-@@W_T\3X
// f\OD)20><:Hc^56#QfGWfQNaU-UD-NK94IE3O0=SaFg?U5+OC)[cB/B<(afef,EO
// 2.QG4=ESIgFWM(C<LC+\9;BJ+4LZ-=2NMdJdcbJ;RT?F(K-B.(Rf9Z=DC/AV&;W@
// LO)UY-a+QTXICb,I:0PIN[1dH79[GgT(47<,gZ>2=,[-]d\A^X7;g6,UC(BZ.+:2
// DP^8?(6_b#afGKC.aVHKN+cK)SK]UZM;2()_VCEDK,C_JEI3^-@.Y>Ua<Bg>0&_@
// VQ,U.G58:SD5RL:ST=cY5[<7Ea8DgLJ>e\/CLFI_6ZLV<,^?74AY:a3M8?fNX(UK
// TKBFUVK5KOR+MeTeMKG\\E/_]VXK(1WZS6M>,cTc>Z:Y6S-a(W?5N7&2;MR>Ra-d
// ,+6[Vb,JS@UbSV--G#FO?2<:<1K0aB&Q2f3]41P\G-:4Y/WCL&FA?2-YSB=Oa2UN
// dI@Q7f+=AWD>=PU)T>GA26^G@TXM?Y-d^1Wd\HNFY)b)/WggQ]<VD:a-/^:8YE;@
// a7PYJ@dIb=2-HLaHg9F?242bZ\S.N<QTF/SYMBQ^Og?UP5W,-Y^4UHV8;LL8#(N@
// 73/&C;A_I/:4[[[>cRJAQPd+IX941->)bW/RQ-LVH:G/XK<A13f/.X.TB)LX:YD3
// ^?U\Ce6B4P::3Z2Y2Cb67HgRNa7;B[@@Zg_B7BU<c9eHQ/3af4)L6==9d?<2-SL?
// =V+5TJ,dXZLKa,/QcSE4,JAgNLcV#<-ZBbR[C8LSO?HHNRARc3FKF3),47VcfJ^&
// #.1?2,;+XAIZ49L.>WLI?&9.-Td[I^HdZ+0fG[PJ<ON=]@I4H[fI#J_L\N.Te7U9
// +8]#bQ]\fDb>bd0[/6_\G^GX,(<\F;@f.D6W9MDB\UH&T?fVPSY(D7(cF9^UdRCe
// ?Q>B@V@?,H39Z?5)@]O5c2Z8@#G?KN;A@8^<)L&(M?TXCS0&+gOR=R;Q^-C,S7+Z
// /T)50QU_^\EeV;cC@YJTc@@&[0MbW/K)MNVb+_eA[G4YJ,54KN.a4_cK[YM?L3W@
// 9N8)d^d+b>?/[ea\S7=8P&GUI-2gI)_)+:#.G/8[gVFcN08-HFSZ3+W0^b;eS>N:
// ^M7AP=TaJg-&PPcgSIcJ-5.2+)RKGX,OaG)V4)W>WCJaY;Zf]dHRS4N64P1;=+I1
// LEYJ^^.g7XcSe=B]4gN#c(_:S#F<ATH<6\D1ZWO^^T,6FDQ]Fg<I<PYPNCc\4E7^
// RK&YQ[DV^264S1JPWcMYA]eX#9_AIfB\7a[:B@\<f1BI];A0C_dQ,;gWSMB8aJ:.
// >W;b8SSX60a==,EHU=T(&-UO;U15CK)6]5P<BMPZ#B5[Rc6)0R1&+,Y.VGB=E[1f
// F50#RFX2-CfZa3QZ+J5CS@@FU/EG>f)f@>&>9@]CYB=7UdFB[G]&K>D@f\AT#R(#
// 6S6Bg+IYa,A]XODJ4E024YV3@9KfS?Q+R3\d5eNQ9^#TLeE0\PF\@ACBVQ>3eHBV
// )[5VSR=LgV[YGC.=-:RD^]0L(&<F9Z21^]KFe9ce+dN;=E-A1-AGIZae^XM68/0H
// +P^O).I.<&[3RJ_SPJOTH7=Ne(O7<+:@;Q3f:C5_[M5,>&B[-P4ATT&@SBT\#e0M
// FeWZ@ZS?4HE_HV;YRgX#8MM;HMLKg2aH:PNL.Za7/+@SH>]g#KFN=_bG82Z2HeeE
// FV.#_MZ&^83<]#PIWP+0/?a,@KOJ-@O)?b)TeSHgVXN,D_&I&W6;U+FDI0;3[&GO
// EAdIgbYO5e\dEY)P66V9=C5f\RLcGESY/D1H7M#d7WREK^#IXZ]gf-53EPOaGE24
// DFT=.O2^fFEF?FHUV]+5aU(&]a1N:VRgZ(]?=EB)L[65\X9GE;.7K8#]7;(Rca&T
// ^D.e/LJae=&UOD#?-XC5?.[?5Y^L:AN,3VD>].0\^6f)&<^+f2P8N/^(^TP#-GQ3
// 0M)P4fM?QBIdagC2O3d9B#HeY_4NJR8-@@G/T,F34I+:(2QUFC[F5R64GIAg9D2b
// Ja9ZR?6.O>3@aO3fHH,+)Q5G_eeU?2/0LP9F9R8.gc7C?M2?R>34D.),(L=18e3D
// .:>7TF=cBe\YNCF(V=SHg49GcU.U_@D+@?[LfKE)d&^TQ\9E<R,<6B-@B,24:)BN
// 6\:f->efEG9CXaKTa030b.9]8Mcd;fE+,Q4M0XOK(;;@5a@D0#aY(H1J/A;gQJ96
// 4+N^+3OU(<eZEZB>X_Ee_ffJ[8<+[;:1CSbZa4007gZ)#+(\^;(5>VY#E]@8ACRH
// ^GI7EO_0RDDf/H:2c7STALF)f#CVN>U3+D(g1EBZ8=&H<Q:VeG@TX:KL&/P6P@K:
// 01b,CT#Z4ADXJ3]9>42#,?RMC:&Ce^g<T2_((5AHX/I86,BZPQO>43VAX\cQAIP3
// (gTJG,M?I?<c<4CN28\RIDQf-I/?3TI)X+,ELBL0[Q\U<,QFU:^U#8M&]XI]WLN0
// _7PZcQ]2ED7(OBfV9OYQ3U7/T^+9Nb]:0-#07:_HJ8c@K??PN94^\H5_\gHC:@9,
// M?Q4)JVJ-8eR\NJcLG<)&K;^f(-PK:).>02C_>(.2&(A\6T]K4V0Y8Z&XJN-6(/3
// T=(ZDAIB;[P?6aeKA3/f0#\@J=UIJQGF_=XXX)]+=G>QF3@O1EW9b@IcM)4DH@-d
// a:P^B7:>AS@SGN)&]&<5JT9?ZUIBT56PYM31FR?2L:K6+4g69-;O^7\79c(dQEG?
// QM2,ZZ9^#:O&@[]<6<U^bD0P/H[U]d_B[+<9@_d.aKA1]2_L91+\_#5(Q4SEJ;-T
// eWAJK.A1eE1?#0K9J+,#2^42Zd)=VRT8IDF(T(bFTX5I7T@XJ;QDGC9Td1HZabBJ
// 96M=00J@d(C,#(5<9NbB5OTU8ZC@bf@;=:Y@JC1-SE4OF)JZY_1;;Hcfe5+\1XEZ
// F9C-:GO7(=a@@..^I#SV5[FY\\VRA>#HV<BA:1a2OH0fe;^7=f84(=?g<&4-:eT/
// OWL1SUX#0]&0N,5\?76ge/I2-\-Q<XgP2>Uf_2XHL93cN,b\75(eEfaVN/Bc-f8]
// 2QW[U@W3.O)Hb_KV?-N\-AES<?.f1#49g/D2#O]Rf^@F4B(6eJMH4<&)\7H^/CO4
// b:J[CRVES<Yaae25/L[_9,F]fJ2LX0]B^ed?(3B&K,]_ISe:\+:WHaSC8#dcFbS?
// (&@;A(<,(JFP&Ta2K4f?7T/I<]/PbfZT5]3B19b[26,ZAQJ30X+@M_9IfCAMAJcD
// -9(bECS+<4c(FR)=1a?I#F0c]W\=_=TTFaOY]^4_3Y<O+7)R1N8SJdTDeJR78XZb
// <b1H8^CE/6MP8X<fJS@b.gI+e_aRE?)H>23&](3HG@H^,L1+KGMb<3AW_SQR<OQg
// R&>GfN7M1VL2KXdQ//&6)7<JXUKK\VWRAdcFC#Y9WF#&\:\]WVK9>GZ,N-e9@Xa(
// W[+8DOgDR6RgLQIA0D38V4SGYOE-J(J>,BOE2c6/+B>2L+YQ>K)0?7KLI(C^3FJY
// 84R\Ag96[F6+?-RO/(88LR+UeY_Ya^[-U_cT/0&1+4@8YYHgL\#L,.52.dFfd7N9
// +EISBF:92gIU1d8(CHfH3G>S38d7V\_](0E,-A7ed?2[+\\g)3_G#/d8)7NBHZ\Y
// )0Ce&]Y;F9#F-+9/QgU2DY,V@R5M4P;]/EJZQPN]OAdDK)1KG1^+6PgG&8(^^Q1b
// @L)Z1gPQYDAd4>B6-E#A<I6OL^GR=7bM-DGQVdB1Ye968aQ6BLN7]-=HQ5X[eHFN
// R-RH_21]2UK.+fEBbg#Sb;HS?[9cQK)a3S,.-QIWTb1\2,I&N/<:4SJI,H6I<.#:
// ZN<0QB36D+M7YAUfL#<DUO9>&.WD/A?2?3E2g#T-<37g](CWZN6+3V^Nd9ac0K[J
// PH3.a\K8803:)=R8DB__Pb#PfUGHZSCJ5e,4:SeG18a.PBPP;^Bg?\9c?/KXf<@5
// T+M[_<AdQ@PaLb).+]7NBdB==d3dYc?(XH1<31:[CT(H63ITE2bRS=N;f4?cQ_cP
// FYeWbX[0M>90N<L^OA0)3S>IC_#.^_d\W&0a20>W)B;WRR4N5IXF;EA@Y_/UE<A1
// 3H&X35=NT;eF;Md49bg:AS]28^Qf#=C?7.93D;f^^5Y-Md9_g0,.X6=RU3G46DTI
// dd,DK^7/A;.Ceb_5K#AV>a.Q.IMN4??0=C06eISbABGdTSC<aA9W[<0b9]<6CR?<
// L7;/X21bd.0KX,IR[6ZIBH:Kg=0V9K:1/M8S>5Kb2\A2>1fG8f:,09-)L28T#B:Z
// ?)7W(8Z=-Eb07NQR?6-BB]W\;9T\T8O2QgD0QVD4_8d^9VF<0)<K@592.9L&T/P/
// :)Z8&3IIK6bbO=#2(.\T_.O,DdcP,=^K#dGFRK\-X15OTH(,:[WY=4@AgII_09:8
// fBN:=@^9WbH+J(e;?ZAO.M^baFI<9]JFO?YTR.G@>KG)gX89+TFQ6F-,Rb\=Wf_2
// /:^(@RZe5_Q9RVAQ8g&==[70V>S:EVb<:?L@]+7D0.KEaXVgUXd(XYdY1TC[KE5U
// D72SC#;b9QZXA]ZZ[V(I-]<YCLeR6I@S9NV>IIWLS:9BLF2J.FSI=L7TcK,Y&&]<
// B,&MWeGZZe-\XFc5e9\J3/Z2?f@))Se#eLJWMVO=9f]L8/TC\Z/0;UZDWK/fXHMW
// L>,SGZ2)BceMfD.<afOdC8CQ[HNH.TFNgRRCH._Q)/Y369,S<63AU#4d+1TZAD)6
// ?VW;cZG?GHVC^#e&53U\X7,bQ9eHOVN+:Y;R[7AV8cC;@CY7GO0ZBD=d7QdMJK4M
// Sc_N_gN5bU>HZIYAS;:MH+,]Y[PYKb;8<40^Xg(@MHX2<UNK=Q0E=6M)J3?LGLe0
// d(RLDRK5:TLH/L+e\b9P>T)KFaU93fJW6WB:_@98<KNaKIGXOEV^@5(UDQSD61-L
// B0LegNe4A>HTTFXc,c46g,9EWH\M,M7^XDIAM<L79RZ?5J)G.\>9gE)B3JL;C-Q:
// ,HW./YUdZ8F?X82Q.;7J+^]I:W8-4U743:&>@C3#Q=a7Z/VMa<A1SafGEWK3fcdI
// 6EcM)3D5-Z&^?O=6-WC++[T\[+4V>[1P:8.#BC5.XW5=@Z33WT_7B0Hg.X>cI4<Q
// gZ8Wd^McB1F.D^>B^dBH(@EPUUZ)GF<XDc8=YZKdKKT,_PJ1GLZ]C)M>?[&K:&-@
// D#UCXLff)61E:bY8SPH,dc>ZDcVFM@@3@g>C(T8SZ&IU<O>7FTcPD&3WT/RFd1TX
// GFFV=BS=DL).c8><0W;.Y00DBcLZ<Z5\1&V4OV7NXXA9Qe+.cZ9&X57gY9bg=\K^
// D.5ZZ..D=UV\1eVL348dGd84?DIN]eNF+dR_/GOQ6F053PJeRO?C9W[GfUR,R=S5
// (T[HV<)D\#Q#&KP9<8]0QSL5c89Zd;V(PY2d[SP5fJ#,\M;^GW&Ged,W>N8W(BD/
// S\\#fKKMGAFR5H6^6fH_IDC.7Z.L^ZV76#TL:U(/-@6-ILBaS9e^IQH[BA:EQD5;
// L+,.Q.,>+=O?WS9P.4KNXdd_#+JNcBVLJ6^N1&M3_IEXV^>>[a\c0BTC^>,;8[SS
// dVD@+Ad(5V1@9+8^S+(c<VcP(9c_:/86<J8@5\&72++^8dH0GaddZI+GDT;a>HW7
// THRN07O\_.eMTI16fCE)9.Hc=#9:_@eK,HR1,ec0B/6X@8)=gW:MNd307C_2d;+f
// :M3SZT><e\;=G,-G0(7>COJ:GLW>O1g)bUK#IgaG5PO(#JJ5Y9[UaUBHG6W<<KVD
// (BRDB1<BQTcI;MfaSe3>_>4)G^FEQ\dOU&OODgA>R_A5ZZW/Y,?d&E4/S6QV(T+Z
// 5H(\)UNJeAF70?QH<I.50AY^:4bf-Y5QDJJ[0W2E>)dZEc+g^cV2?8XbV3WXf,+F
// 5L.GMP\.egG]3Q1L_=9^,f7<Qc()ZL4IXZ-APO@J\LJ5K/1fZIgeN)P9NELfNT:P
// =JRTPM6(gX5C0@T5;:R/NdCUK7_9bIe4_)c&@4=#]4IJ5.;bf&WW2fWa1N/_LT1=
// JU2X\WN2/Z<5C._.WILLO1]?JeYU6W?LFGD6Of-XT^g)\Z[ae)8C)#VVMW&6H@Ef
// ZaQZ-21ZWMAD9V(bDd0[?))AH)U)AgXM=;Af@H;F2e#LV.1VdNX/K1H@c4F>+\Ge
// ZTIEM[@95;S)b[KRa#IVPSVT?Q8;O-2HT.dKF]B)5?U\V<YQHAM0\+U,BF_Kg&cb
// AJ]UdW0^_U-4<.](>VYMM.(\0U+B#_-#T@BCP.1G71EBD.[KE0eDg=gQ:5(Lc4/)
// 7L;5f@DFcW2dJY]0T19MfGSH_g/E=DDI#b3KW+bC]Dad1AIOeXgdDd]9?K_g@6Z&
// 31BeSQPRbAXWM,CE57-7I4E]SS(ZJIQ)(N7,):_f[e?(gDgA\Z+Y-[/-+,DM-5X5
// a4N2_F^[d0-Zc4;7XbC7_BU6RU7O.eUCP)+_QJ/>-7Y=#(1<+-^I<a7A)ZXPKe(5
// (?HC\-+g>0FNIa&67>QP7Kb4BX#LfH^?F<dK[.TgIGM\H-CcfZ_;K6\[71JMID@]
// D&G+[L#-\BU\<3S3TR<CDO;5\I#=Ig=LfTYRUD_QgD.7U;<O9NKe()Q#OB:VRUI?
// .>E_-I(g6BQ2WWT\?/bFE9A\QO-4TRLRWb)O?WJ<88LDeReJF>\F614Q/PP@D>GH
// 6Y(F.UXD;@5gC/K)[UC71Z=9#A5P_R/.XOS2F6X)gB3bQ7[+YUNeV3>O3?/[L,0+
// AE_,W@3f)^JVKW2B72E]39:@5f=KT6679+gFfEV=Y#UG,^P94Eb26MQ7bT-((AMD
// UNcb#d75\8K4e-@8F,WWK?Oa.M2M0?6A:DAAEFCHJR7?,HM3:8Q9G,;(GUG&KE.d
// M8@@R50B2<S3O#?BgY@#P(87XU8g0T?B7g#ICe9RbIBYfXN@5Z4T@(<3b>)6[9<U
// ]_.D:H1<8N(PIO[VB0SAOA/2SeF_-dZg65g1&N/(QOc9LUO4Ta41[#IVS<L9LZG&
// (3]0]?/HaB>Y&Q3V38Sc=/JE]_MM/gcA6E0BKg]IC;->T5O)cXEgcd]8FM^1;;Z;
// =KR4)K;X^@aa/W:[@9^7.=56D>35HUSSE.d3T&JR<b]-=4:dLH;G<^UBg,TVdaBI
// fd^0MIW_9)O3A\D,OT[?GC4BV#e=g_16IZB]H?PZNJbCOI=(-7Ze7,<SE:<RSTd7
// M;_;#5^7P@bTc5b,dABaXcb#YD8Y7be&.XRg<(J@4ON\dW7]eD/_dM/6\QMdO_>X
// MY\:dX0LG2^6a/(?T)ZNPgD=If@2J2JN]+&,I@c93c>Tf\[:3YMCZO^\50L#TGU#
// (26BTP;M/3?5H)U=[3_=aVJ:MD.&2aE^UbNa:;W)REKG\#>\@[)JU0W>,c5J5-1P
// ^V)F7:cG^bKcaWMeA]dV7N#56ZPZ+0>\[WN6<F8953faG-LELKUL;ZbeA#.A@.;C
// 7cXM5QT]@Q0TH26BW?<fVV]EUY/1a=ZaH=f)c>eTgT2]BX8^ZG2^5/P?AIHVFENa
// ,0P:DaP@VL6-V<^9@E;f56S0,RL>fF]Rd3PYPa1Ha:8eU+/10.O0)gH/-M7B1==C
// 9A6Y.@\-GNP/;L1A&ZFC>H:]^ZYS=+9;bV:WN.&>PA)U4-4:,@MGag(eQ1AD?_&]
// 8S.B=W=&G\8I2S/5,)2Y4KS=L7&F7dBSH0fF(COEgE<b)e.&HR-R@=\&P=TLd@MA
// \_QW9ID(CVAGE7,VJ16M=V82N?=R-0EZRT>OE5B/33W_CQa62X6Q+\6fWdCSNN<B
// ]RdFACF00BeZI)0O,EdHg#E)A-+7_F/C34=NVcg2^,g[VY8WdL:)4XS8&dM)VP>_
// XA,Ba<e[KY,\eA55<Z#N;If:O5#7_QXDdG#=HgYKF7d<A9.#88Gb9J/T\ZVEcW46
// ?&CZcS>LNTP.12>gHC[J<N8B_#/ZHLG6S9eCC8LQ1=KaZP<=J<P7eP_gaL?/PBc-
// ^@]DX.Y:eG3XMEQVcPQ<GS@M0c>J3QQ?48\R8K0O-;agf.(1_gdLR6KcP5M;F;g8
// O^BE_-6;;;Y@QaHb6<71[6ZcN(c]IK+Q9RL#+WfY=#f?>F\\gg[G>?>_LIgFYd,[
// _HA5aKJEOZ0dgBIdY086]PL^(:\4V3g#\]&ZT1=b36_6K5>_G)(IT;#MX07QZXe4
// CD4GbUDc@1\I3>OfI=QT/6CT9a:OOLTXd7.bQLKf6(3[d(A[d9aS?a]C[89U+TFb
// 9f&fLFDK1[H^@9EOFU4aOeA##8F;:(R4e+]<^.=gW9WfR:a/,T08Cfaed+?7_E64
// VeM=MUgGeG96S.fCa;Ng(M#f9Tb(>Y=1K]8M(;B4ELF@?+DW>Z&T@T/9X+f8_L)Q
// 9F7[e=N.S.L=DQNU\B?a=SBdc8O-9[WMXKTXM@aZQS+=MD>Pe]T\P_.7]L0QTZAO
// BN4afXHHQ[5P8NGKR?fH@RIU1RJZb+8>)S+?5/E4W0;JP?YOa.R04O@XAHE;,/G:
// XER<e;7bSfQG]G^8Le_bdXD8XD1Z6_:@S06]K7f=8P1P@4_:-,=1XU8PH1Z;&??+
// d+YA-dX;Qda/EKMWKJ)V_ZC6H#QLcM7KDN4XeeOf[6Db7,aE1+#b@C2_EBaKDbZ:
// 2[3S)V^3)V<Z7IUPa2(,4-.\_Hd^S]Le7C-4=Y?P(,KOTVFETD26]\_]FL;SO;eZ
// 6>O9][R?A5P[ZJ4AJX7+82YF=3MB,T+cYLH?:0I_W]>+1J?Y]X4;,cCTV+;JW2gP
// 4VTD5)c,2bCb1^F]77PLQ)]@S9+KIXS_<=+-+>0&fZ)9fc[_BF5J919Z#1K2DAAB
// 41@J2=J=P/I0c]6edFFD#QS/#U;KCU4]KVH2]KZ?ZS?2LF<S:I6+cO4LACYA[?RP
// 1E=AG,2?W,I4=I1SbAZ),#Tf)SD.]TZ@D3EeSOET6V;_JB3_X(R(K4Q-;LW215/d
// X=85ZBWCJc+f39#90bV#E.T^_M))4;HQQWS_5bEOIV(cfK6?5GD<F,?dWd#)+/If
// +307T^/;9+,X_SV/53bURFe>&/9C;Z@9NR::-;(Ub1_d\)A2<:^2Ic>@<45J->77
// &DY&U(SEZaGU2F7X&B^M&SZ))@NB,\Y3[?JU8eN&Y_cQ+RV4_SVECfaOK,\3/-4Y
// JTG_))HV<fVg<6YTH;>XJ+-9E_DK\0BLZ(\;^#\CcQdB&[]AeS^WA<+DF#25GAEG
// Q4cZeBBLNEa.-e,]+cAW-<acX7ZG+9_YGY<W)(W-:S?.;>PJg2Y1XM#H?aVFEfG#
// R&>f:^ZUBARa=0KP_3YF=;8WQGSV5b9&&4=dE+88fLTZ@_[:PM=7FQNC[E9XVZQc
// _aT^?BUMfL>\F6;NM]YcNP]L2/AV-(2?;O2>99M=/3_J9PU8=eT(O])U@6P7]:;T
// ?ecQ_1U??228,@Z;]#DaA-B&L0C\SM@XE,9^R,>\NLM>P,/B-OdJQ=KM3b.#Z)9@
// 2BV)BT<Ec)J^cMX1674IG/H,S]4g/(B/^IF:N@YHGMf@ES=BN(T^aGOGe7Z4c<A0
// S\=S353KFF]<TEd6GQ?O/SB\U7K46)XRVE;:@[YO1LW/Sg15/6XU\]3_,CL(D:?a
// =>8S?4dCA:)6,g.;aE1(cEF73,9b#C>J5L6<K3Lf@R0[b?Q9_/ePRCe7#FF&bId9
// DBQf+N+3^7X;:6IMb1e.FDK9OBIK8<fO0:g(QJN#2<Pa7UZOF/RU&3=P877IC2O_
// #?K/bcYffOR=MfUS>]7TfKI@-RcVDAHaWVZ^g1KMT59P[fAG1+XJ;#WL\(S,.dD@
// DCLX:M(g2^5:6F3cIX82/J3)&11VCP@b49J]7eP[F-6>HF9+[\_Y-d>_aT]1O)6W
// 9Y_WVQCa;[YKV=d;ccK@;K()5&R[YG([4QLNC.H9#B4&fPU&-[F#5&(5BL<a\eXE
// ])XbE:3Y?[=H3CGRRQc+H4N>eM?:RX7/S^:4W60.OTJH1/]Z.OF]N4/P?eadeR10
// 7KYKVY-2dN)\FRf9a]e3B#=eBgCRAJb\^V+D-0UFYQRYP?,>8-H)VJU#3RY]c7&2
// JWK//+2>XRZZ-)/bW^VVF@aTD>.eVDX)?NSW6-TaUM&B5f3YEId0?b<ADB9OV>0_
// fL)>@cCXBTH?//7D=I\ZQ0@GD_UK)#FFQ=5H.:K#,=A:1/+M,.a>[_1\+ZHYga[M
// =77B9(g+4)WP/gNd2NG6E=_.&YU0PYT@@0T,BCL4^XHP)J5TD5,UgWd1JIU#F>#W
// E19F4Af8?Mf8+_,M&_8J-8OLOCX3QA=5&9G,c)^bfgO9WOV[(@_[X>6[Z02V5>c[
// 9#)<?983b]/LSe5P320(L5UW58BEC)6N#@gO2=O/J@Y/JW8GR_:0Q;,S#7QK1Bd:
// WVD7X#HY?be(:;:DSbUdaR8_H1BX&]8>T;gN0Y-JZSd9W_MDEQR-T&KN_WCc^1S8
// af^c>>ILgI20(e8=<2,L]^?e>?PfAOVQ1F+3ANdO)#@:)2/Zb&cX_X;1P\_PLTQf
// ;3/17CT[Gg3[\gg_Tb4=#_255.VWZXC\eTV5gM6eg[<D)CcK5fVg:VTCPC0F-V2F
// c)eG7df#I6:(Y)>9[&.,?P]MO[X=\X39-;+X)R^JK3NIID<:_I1?[[O1?EMN)ZTU
// KMXT6;P[FH;aBgaTR)WT5Q/V@Z0U3QA/YNXGfNVN+CeX4D)_3:S5J(VTR4-J,@^.
// S#)<,?OZ9]/HNEfU\5#A8&^>W\gGQ9W<.IB9Yf_[43FZ:LEJ+LFcX;9V9MQDDT&R
// BJ4=?K=bIZAWA639MZ2U>^/df#Q53JBB5a:f;/b6OAfC#D[f7<Y5HY@NU+;_5-/M
// W7c9QXJ4O];#f#<(Q@J_.4IDY?QFd&#Y8\\\(@[_ELJS+WD_<R1ggDT[f4X5.S<S
// 1-9eW>E1VKLO<_IG7a#)MO(FQ:AN;O5bZJTL4O2WYce1AP)FMV[H-9NMEfaN@/D6
// :BD&g<95B?\H-)VLY_O+;(?=Y(#M+>7J:8=e3YTL6OY^K_1T56OY[Td-+PAbNa1U
// ;E653>=FTg1YCP;JJg.\U76VCdeXGTXDI;6ET<@OQ=>?QKTJZaG0A7+B>>f72G4e
// 6R@[G94eBE8[G_FOJ>VR46K+BeE;P5cP0;9.QFXPRZH]C[D3#;@^_Z,c[R(HJIO/
// J/e0QQPEZ+)63>69H[0HDTGcOW<V4=.Z\,VLQgN_Gc+OST,(Y/_bIP::.g,[a)8e
// 2HA<#Y)J-L3QSS-@K-VVUDcG777>LZ@YO&C7O=+LP6[0)RX4U_/M..9-?CJ\&WBJ
// IQ^+Cb(5ZE9J/(0c9UJ#:9N1U[#&cDSKcV^eO)[/:76Y[Z9Nb\KQDGXM_;#,f&SB
// Jb;dQV7Y.J\<3YI--#^D3R0=]YU0F]F[I17Y0Z^:RVR.8BA0MO3D<,H8Z3c@&0=T
// ;fQQ44V\:-JUd(K\UF4cGW.7W/838fZ\#Y(3DM(7/.)UHf>_#RSa;d0dO41P>Kg-
// V+/b0AAA-@G4,6Z=b]A94QHN;FLRB?HOV9TL,XC:HXH5K5,ZW9e,Q,=-.Kf7Re^,
// 0ZAcLCOFM78#+5eW&([3TZH78L3?KK.[?e#Hg8a>/:G6W1U5eg.RgbcU7/?P7E7Z
// -RM=U>gHP)dN/JLSZ=7Rc1N=UD=T=R6TBHGJBLLSZg=/VW8BR4O+WZ#A]D7XMNG@
// KD:E?L,.7f/g_d<2aeJN?^GH;aEg/b9K+L,=VRY>BDgFAH<6S+c[6<WNF,IL6BR,
// #&f_d\I?F,NBA4W7:fRKDD5b5dC^S@Y<.3S4F&3D35NR+-a2d)Mf9SZPF@]JgaCL
// 5I]]4IY+N+g&N7DS]O6B;1H1H;]NKa59LC[R]/4D9#;cAX-(HGEKH?@SY1I\46FM
// ?D&/7cDC,L7MCHF9XeOe@fJ;)aN[I2=H\ZXOgeXNfE_b[0D.]2QdHe[WY081bF&V
// AQAQGPU.)I\:7RAS/>f6R?<,33]L_JZbLMf)BS2L&T2H8.TA-IIW+WZM/T]NbNFS
// 7f&g\0UH+A\_R.dFTT(M9.>?d6PG0gT69faA][ZJ3fC.@VJSH9A+aVbX#[8W:fB@
// gPfe9W\\g[A1X8.YQ8a_U3WQ>:)@V7\2PEI1fBC4_&WX,#=.ZWRYMd042;\=NYHJ
// #LdW+:67WBNN1dD70_HN2Z>)H[4UT&7GQd?Ad717@0)(V]YEe#TZB#KJ5OK&)>Y;
// AE3(gG8>/M_IIZ?VH2bK3[UgdBF#d0_W^#_W4ecGgTHI;6b//]N-SB;Z,PZeEc)7
// R(=9H]8_4K52KS67/_Q-:?_CgL</BES?VC1^<N@S8+]Q.ZHUA<V8b?UFOagZ?Ua^
// FUfQBS0F6Vd.M:/9@:Nc23<T_K-CY@2fOe8UbUH4Eg=@@AHZ@FgAKd2AD>f7^AO6
// a)^P7J]QLM3/YIgKJE@(b5(/D\R&EJEGcI84RF;ObTCgIMG#a>UPF2Y6><cOH&8N
// N]a5)MYW\9RVF\c3(Yb9d4LGB92TXT-Xc5Z95DQVZ-G/ZXQ4K:UC(7a;JgMD]a-Q
// Y^H/>&L>S[ULY\Y,T&0U;2)L>fdB3XJH??)>ddf1Y3<CGH/Yg;73DVBC3d]:7AHU
// V.EKGZN##&#-aW?S@;fZWP?SWV^J2\PN)H(J@@d7<+)2ZA7J45S^U:,#H1+.TNYH
// S5_dAJ4Xf9B=>,\5PS@M;HJg;c1Bbdb#g8EE:^8^@E29@JX^PLRFY<bfR&U4LEO&
// .G17c9OB:+FP7QaHSW5FCf9I6?:>ZLc0>g:?ZccG88f-BNYVZ5,KOF-:M7B3B>J9
// [@ae)FUBU-X+,e>),6L.4U;A+K0@@ObPW0@R&NEC9T2Y=,:QX(L55f8L,La1#S:3
// AU-QT:^K3E@9gg;7D2R/V>UIP^A;+c-b<SO&=+[_<F(N\3#]2CfZ;Z9Lc-AZ,^1_
// @/A1)K#geN2&U6dR]W(?+_ZB64;A(c+IDSdf1E4>;g0##bc:0K_(Y^59B,[d]B80
// VBg09fJ5&)gZ)>E]=Hc.S;BOC<Z/WHYCG9VD_5FMN8=]@+g,:X\=7_2<+Zd11e-A
// YEZ>RdF\O9ADI=g1VR6f3MK:\5JMc+3-OPI(8(f3-I(E3IK_/13a68GY-cP?@;87
// 2_,KVLKVZDc@c#62[AMOJ6)@[.-0S_8a<:SB],f/+D+[-PYUQ;L^2/-HVT&U@RZf
// 4=M87Z?LB1RB&:T2#?/K=G/V>\C\;cJ9B3@2=3EPVb17<)SWHLE6\CT+NC=FDJ42
// M\PSB2Z[>:;5adTKIeEE.F\:EF_Y5SaZ^Oa&^:[7a.VC0;0VKGce+6;AO5R?f433
// 3S+A?aCF=bSR?J^QQ0V.Z<1P.S->9STBEAA:^17De;_5A(G6b5@eDAdW<O_Z=gG@
// ]Wb?67XQ>N&7.BHa12OO7?19=T<TM]HGZ3L9+P2BFDbTT,0F#bY21<_2CM=I#D:a
// #B^Be</d>_\A-GHEd98Gc60=_OgC:WD+JZ8S=NEKP1HF78L@IaaEKO)=U9P_=_;(
// gScM?RUf6Zg&-5aLOY0#\)D<1U8/KMV6>f>.OKJgZ>G([d@e4H\_F3A2U5I82B<e
// fJ1fAcYMJZW#1)[?RQCXZYFC\1H4D^4A&HfT5NI(^5]bZ^D+IA1gB\G]aU@WM-eV
// USE=+,0W[YH,[Nff[65c9,J9d8d=P#63<g_E/fbDC93K3C/PX(LN@.b,]8H+]/>I
// F-=D>J/WY@P^#ZO>f;<#7D(NC.2@H?1eded5N<b)9@U7b0,>Cd/2[a+OV.>:2f52
// 3gdBU-GG-,S7gKf=CY_16,1g0EJ8W7e94c7<14XaT7]HL8T^#TS6ae>)>@..@Q[G
// 0O)GQZQ&[4:3]BZ&AG6BgK[X(c(582T)6Nf8X]6D8-T?:@4Z2,_[2gAa]SRK\aaL
// f#^6O63FCH3(UY,TT@9ea>@:HJSdc8<].VSLP9LJ05U5<112MI-W0,Ld:aV=HK3I
// [-&ZBH[6BV^ROW8GcRFAZC\Z/UNXc_NI]3/bR/P(FUQH<Z]K2aP31E;f@M?,T_B^
// d>8-CZELPRRFHOH>g\M<50Q0F85ZPAX6>IbE&INB0eD28IbH.Q5(BQG\U[5)-C@5
// Z+Z3@Ba=#(_=C@HX?MXda4M<ZKSNe\<5OS)EY8J]dZYADN&Jfa&-;243I<=FY#L3
// c@+beHXJ)1LU>06\DdY-5a/bI^\Ec7J]1F@79Z@XLL7J(<8F2+gJ]He(Je-M+d^Y
// F=V63ZTBASTgcFTdTBK^E8YbA^.cE7B46,EOXYGU364g>VNM1.CG2HeD>ZP_LfX_
// VCH+R<-\8(&QB?N]-KF9IS(A7cbgV)7/Q\IT[K7dLN<E5+0#/+Kg_de3?N--6DaZ
// b9VXg=5=R&YEB(VRe?KOT7@Y&:=)35QVANN90KP#_YBV7K;3:Ld5acd[3U/;5+AV
// 7W+:9.;9a<7c(FLFVQMZHZN&X;@DdF/V)LJY;d9=PBNFcaLK[D+>C<RXK6E-.Z[E
// ga^1ME\3NVKLYNP/2:f7AFS,#:7,=RTc2HfC=\<KKD..c)FEBdD,5EKW;.X5ef0a
// K);B<:U51XNWNX2a0LLfG(ZIR3BL.B\STEQ/EYS;R7[]^E87-TG9UA:G:8EB/#)9
// #g;05Mb5W,Fc3]&aW:IfW-D0FT=YXX#&9=(\[ZOM_dPH/W)R8ZRW.?;?Ta;RZK/)
// N4N5agD#D>07#M\B#85c3U1#\ZFP&PBb1IG_+gb(2^3D-f^18+#>HQeQeg#I9F/,
// FV[.MbPQ7(-L)<<?G6[S/78^;a9^Q&U30K,R+PSbD8S(Z&]YZ/^f^>H]@_<;GB_/
// IJfeW730.83#G+d^M[.HBE6=7#3)6TW,92W^@1SC@7<RaUd7-SUX4+L\XbdgDDO5
// 0JY7HE?MIO,\E=d<>.,BRH-6WR#_7[KB43_Ga+cJaE1gR3^g&=[[=EV/366ac)cF
// >UPU8)</XS9^eOI7^fO;0BTMQ>a;PXF.+E+.;60.b?@1-.]@C&AUM(5BgPDf@.Rg
// SF?(P6E&46UOP?>4GKGg9LRJZ:;3:N@g4Z\8cK<T::Z>-V96:83Q?L7+@^[X\U=d
// \<1N5eX=M2D,Y(D6O:YZ0gb,UZC:FaSH1N26_4_9Tf>84/H8TF?S#6UV&+2?M86_
// /Q\777<f-+I>.6/c01PL:]#ID(_7)Gg2(;AGc]D@0ABHWbQ3V?Od\1W/D/Y9+@:H
// G@3-<@V8(11__\_UM0_LGB\:W/VXBBd)EX+[c,7D5X<-:(e?&;#[OIbCBLGUZC<9
// =8/Y)U0AdO\P->bOCIZ[4c80Aa;XQFJ[D&f^;,/7DI1-ZPHfg-TgeXD1??9aN(UV
// +\3A,?ETK.X7(4gG47KOe3SF>81,2\fVB=I,OAQDQ94+-]gD.?1=\/.I1-8fZI&e
// RW59gOWT_;5P5Y:),RVGQ7ECFG<8;37a2.QSE#a+S>]FI&4(5c_Ia;BaD2E;I1J1
// ?8>65+2;\cc(Q/bd<=:Y</5A05&&1?b+:I\X+#_V:8,HX_Q9N?,N,Z@_OKDaU)[E
// O4<Ce[Q8d)T]:YO<ELV/LJA>/EE?KP8Mg_=3,\8;c1V0D=UJe[Y2>cF)@A\cSFcE
// #^L.c=KcV4a3WY.I(FGID>K#^.)DcC-)=8ZWENGT?D22JB3:/:SaB0.<LP9.=B@4
// +TRb,59NY,#P>F:0O[.W+Q]<WW+?)5L<gB-=89MGD66;K9/f.ZZbIc^DAOHRcbWA
// NV,S>;+IY)=_IfB>7Z@?@2>YDMK[Qe^LZf87O8-[FTG]+;3:H722[ARX9OT7\9T#
// @F/.>:RHGBR?/\CR@2e1S(Z?RA_Y5]0ZPF0H3,U@+Y>dfDK,P&OV-dBaV@-9>G7Z
// Y+0IR]O:dX=_Ac/;a0?96USaaeE3;)gGcKOc>c@CdgcDcC[cQR[1>5\<58GFXJ&B
// -fQ,4_GNY4fJA74H/d-^Y?)1FMGdU3)T#.L+92,+/ZK[RDR&B17#).]M32aM3e9=
// :+S9>ZK2/\=<L6d^WL-J<WWM]OYQ.DUJ5?bN=bRg-9B-#<L2=bMYJ5C9<W4VMN&3
// ZYUc&^P@H+g(JGcOf4B,\g@(B(<7W&RRd)[=fA=;]0^e(N;9\<;=,5E6CQC&VPdY
// UU\I5d@KJ9JZ:Y.C9JX\92<A_EF9CEH2VTS2AS4E2>?B>PbG^OM(8]B@<bIa&=Q8
// #2).&2,bE5:L^#6543I)#_E@O81O;TfbKKTRHHPCXH8+PJ\<-<KQc086C\c7Zd\-
// &-DPPH3f;5SA0Wa5@+3(P\eGSaJ3\LbI]Y^:F4A\UT/4K<J@gAL5Z1,WPRPAfNa=
// [(^PJ>?@7JaE=f=)FS#EdH9[M<WJ[O,B)]QHK,8WW(YMcYOfI,GWSacFB4YB&1+O
// YDPF@9.3Pg_G]4Ac5BgF(I5]T,)>/+6)=3ee[^DBb@:BV_W6bH>Y-XQE#)CSUAJe
// _6B9G2)?<@X9G(14f25JK)[,-9HRWAZD6LgGX,#0[4cVdI2bY<S&J^6?9ACS-+.Y
// S1>BRRG#H05-e((D:44e64UOFgN62AFL\]FgSD_(J/QJ.][\ANK5.fUZd2eB&&:N
// a(MBW;IP5<TV+1?6[-<<_2TDS,9/9U#ZR(LDJbf5G2Cea0GNZ\c#JBHU#0214^#F
// =ICS[K+dg:EFUW&6ICd(20_dV0S+LT52=C>R\NFI/aJf\0+#<O[&<GH9[38e-g[N
// &\;:,:V<MOcAb,(\HAK.LMN8//BKE[T^.D3U).5Dab<H&9:4Z[Q=Z\6#bQ<4]46^
// @;5/3=E_=f2/FJ8Pg).@:b4M5Efe/3MKNDdWP.(S;,A_>@4<OC9?1d>;&;V:g_B=
// _YS13U6f0<Q0>CP5(.DWL11DfT\;QFf_3E@_AZ&08-aU2@a74=1(H/)37Jc,:7I@
// g@M:Q:2ZQYEf:O[P#DLc60;N2UgR03Z;NggJUB98_&T]#X3I5U6M/YEC;<I_S1?6
// VP5VP1F9(,+CQ)H&IYCJYK=E@7VL45RGIG_aO&g/[f^c_KMQ:]2FfUMgK1EEEUP.
// 4,]._D0S(C@^FM_c(4#.4aW6ZW&8[:8[6@Dbf,fUPDGP&U8_\5:J6A3JS752RAf/
// PQXNIZd-O,7T>4f6/,\)418-UF:ASR&gNW+\#aU6DWT,3A0>TXgc]>S_A8-TDZFR
// @0c;@0dYDARRZ&JV_<b30g]VN-fe@2F?Y_AUH0;++]H6Q1]5QG5HNNLa0)<)8;+V
// UFL1H7RX6VJFBPST<;DSQQ2A+0BO\:&2b_Z?,0MEV5]dUf3>ebB;^F0eOWX3^Q,F
// 7ZFe8ZGP<<JSB3HNF+KF//\BFAE67@\.R]S<4e_RHY\Q[5YEed1LA&AO)?&^^QdX
// T>KE/6<]R7(9;L9RRddYY\W,JfQN?JN=e<.3)LcHW_?VR-c6ZYD)U03S=\R[M/K&
// <55/Ld4VD8]N;2T)0?^ZZIAVDd_X+BI:>Ube_8Ub^P-<TF<,\HKNH6E(:0-[2a04
// RL9g&TKA95^^ZK/KJ;WX63IJf>#CFAN2VF/dAV_6II7^CaXQW7RNVRE?G\FG[f?B
// [aQK94GPeHVF2#E79:Zd99;bH0E_A6V&f;C#:7,YYBMS2;RB1>RL]g=NS.HaT,)7
// WgC9[QT?7\19]cPX6VHRbL=5>JPVUO;eIXUS[^Zb;.S&LDaI/5_[:YAV/F)6X&8Q
// )B^4\dY3,RKb7ZMJ4(&YE\BFYA4<9Mdc0S\8SZ+\V;@P(8fZ-gO(&Vc/J9&WW?b:
// 2cKdKfbGfEZeIS@d06K:U#&/:/UTEJ5<d^<;(N0^\@2::a0;VGeIH)+E<OFaH6.:
// C5:Fc.9X;5YC8(&@EJc(M.G-0=bA@H7IaDcDM\Qe?-^+)H4C//a1(+gQ^+W)^NA,
// ,9X1KSV9O1YN1(2gNBN4_b/GKd]7W9DV;/<b4X\Z)?^1eV?W/-?8ES<B3XUN5MfO
// .E<?XR-CJ;#VB@8ML3GgBcQPAY@8UFZ06W6Hf5eUCe(\CY:7]bXBgN616&O4,,O4
// U\KC2.VfC^#7fYJ\5S2<#R15gS?2_NC(Q3\^fQM,JbX1=fb.(AJ^/2W>Z+3_4D,H
// 8ZA6=3O+b<c<YJHO/Z9\LM0@\E.;.Db-T0:TcTTT\7X94dc2&945FX=,L,[VPYRD
// bd>K?E?RLXMM8K]a>_3175)6[BKCAIRBMf]dQ/UJZK4>>,<=0[B4NUAS@NPI8F4R
// cE@C3=CCK=BA(MV04ES@g6^_1.S^2g,=\FN]Z_PT4[FAL@A?&&c.OTL):M4T7f54
// 1Y[&McA(.E:g+A+N<T[d77@=90Nb8MAbfOVScP:fX/\1LVBOT61Z]=gE#DN]U=ec
// AOTF]\f&\:#SN/9;^7bXcgYB6Nc4Nf4@YH.gNW1Z84QL^bJ_gE7UGAWDWgP,QV^J
// #;-Qc^c-__Ra7-P;GBA:M,DXU];Wa-eN+5Fg-)31SFZZ<@2Ne@[B?eMX2R9CT#L+
// 8GdF82F[I\]M1=#5)V41W0I:Q3O@D0/-OYY,Y1+PD\7HD@3Z]4Y@/D@JKdEH66IB
// _@8PBL[+..X30aQ=Q1f)77\S]a?M^&A?)KW.MOC@>UJ]S/(:@[<3ZgY>=7=8VO\2
// )][d<5XP8J68V;],SKHY\<cER1L7#DQ9_RDZYbVb:48?(+&?11U_B0eP]U<&(Ic7
// S=]fLK,C4-+F@3McGHJb-5L5PQaH]?WD.]1Lg]+O)eJ59G6)&aB#LN,3SSRKI)Be
// .O.5BN;IAF0dXgQB^W_.HUbX#,Q@=G1CIfSV;:IZb1<2U,;M2=Y?R^^3WI_TMg/2
// N\.<).59>K_A7XDA,K;@M,N)?dBDY2G6eQM^4>C.&TC8<.TS3M[4L,#TY/DFZ&WW
// &(RR0R#V9>I+SMO3?:VN[V?dT^2e_L0F6T,&HM6b+.f4H3Z6YV>TWXd36>/JaECR
// Yg?BF-5NND#@;AMR_f]B2DUL8WX9X>35Cg<L#f4V>(&e];:&L<aW[9?[\\/NIdH-
// (WP[5+FCXWR+-a,SQ->)<\KfZR+Xd9Yb_BXP+&JU(AXVLSC]eK4D9^&HC0R8eT2)
// E;?=cSgEd>//CM2ag+NZA1T=F=)UZNS3C8<3dE30QE0AcUN4d?O9b=EDa,a?##[M
// M4SGQT+#Fc._Y=?R6>[g;EdRKE84H-G[+=6:0d;HRcCRJ#+a3O/KX8_NUO9f^.+>
// P=DQX9E4.4HFI&Y?RT/\#1da3&Be;eCLP4M_6B1<N(U,CE8;.-9E0)[HJXVOaBDb
// JHdV0Y#D5U^R6[ZH^)7MST?/@F5V8Qb;.,Ue>f,];dTF8MeHfde&:OAA6A\b=X?<
// 8(N#eT2b(&N;.9gP2(bIT=>UF_XZ]EaPE9^_,6EH4Ba?gB#VP10]GDa>HI\)a(EZ
// eUd\[7Q)SDZ+#gXEcJRfE/_/RF;XXBePX:XK:ePG)Q?KF1MTZcWL:)Q0R/_.VR&#
// BgC+G-c,-GUI^ZAXNR7>X2B+C1&:cSF1W99Ld=d.SSH4e(Kf3PS@3I?cU31>Ha4J
// 7UCAebL]Wg]eF6HI:UcQ74ZCCD[afW.f>5Y^c#/Y)V(JUDUeQ4I)>d<ZD?/cWDI0
// &RMaQ>S1\-VW)IQNb^/S(QO40GYKbOTI&:#D30@ZEQI3K+b1VZQaWEXb()KV++<S
// AfV6Mg+dCbT>-//cYZ+@,P_2aMRY;-E-N-dO^&.N:\AaMV&+e7&H\OHcM:_?eZ^K
// </87HTF[EgPJ1J++?b1CTH#fSBMV;dL;6GW,/H)>/NM,R(KP[N=F_1JA-6eTf<9T
// ^F+T>NMFaJ.>ca7GeY48OLPHQG(6OXHRLNSHKE?YbZCP#0[X&cAGA@:^+3_/L=\?
// 6,,X<e>)XgVCJga=gD\^8M^M/g(;IJc?g]X2/3J](Nb6S+,<+9?1ZC^,^G:O^8DX
// ?gB3<8f?&26;U:SM>@))4U70ddZMET+K@J2_[H)I),)#cLCD&ZFK7SJe,M@G(]Fa
// J-6#]_?&bC;,d/?QD6c]TM3MYQMQU&[SaZ[+&S[6+HL4,?BSN8I)WI]e:=(V@+XK
// )XGKUJK7I_6RN]Yd8aa5?4HR3[IS6/-A0\IU9>B&a&BG)J(P&<J;-?H]>F5742Qe
// (9P3RTE8cR++9#,1\LV0I_5d,O+_\2<[:4UX6Qfd<IP\;68/VeLOXP6:NE9gBC.R
// DMF)D?Z+bLENBCJV0BQMHK#?JJ_.9J/L4SH3V3a4^75)D5Ce25.>6VF<\.g(T+61
// (5NH7P0eVW?W;\J8N6+3gJW\V#0[<_T;NA/(@>,[d4.F#fHTgM8Re-NbXc;^O)Xc
// S7]<-_2G]=FLA:0:Z<ZZ#:L[]D2e:]+?95\+g<HV?>@S7d8Xd:Re.+e_>fB<FU>L
// 3Pc^VP4L2Z=a?c?7TS+Z5)W\_G\D:?\<aJ.5DN6^&0=<C0;g(7VV2DM9R4C.Y<Sc
// Af]-H9;dR1R6RWd@,GJP>N)8>B=FKSWW@2VGX&4eE^IIfa/9cb>>>&(O9Y[NV2HH
// 830;+9f6CY+1CVUJZVE3ZfZMG27fGL\_fOcaYUDgW)/Kc[@I=U;^MQD5Z<9/Y)V(
// PAN:59GG\J=Y>/3d\6FM,0O@IS+=F(df(-<cG#LRD2/dKPHQ>.M/BeWY7a,Z76S?
// 6C#@?N=AUA;J_PgJX;a7FY,S\WPJ>LA0DMK9D-KA.\44B_7YW&FN@Laf:QR#F\:Y
// 9D64)R&8aIQ8MI@[OI#FLeS@?PU9M2DKE1<?QQL5KCVO21Db&EL(CEO@#\+.4;_8
// Z9);\58g@D55D-=9:FP4(&[aEB:;<c@K@<[I91.-CF)0VDQSUNGI\WW3C9^;0+L.
// aG6=^>G[1>V>S=^bXg</>S)?/Y:6+dTb_/g,KaB2])<RF_5VadT@P>g?bARVVVLH
// -)4F695U.d0fX\bDIgQgA+&I4_[XJL8&S,Ze9fdKS5Ic^&:6Sg2))6XMFa7Ab=V^
// O#d1^e)JQV1;?SCFJ]NM.6YVBfNT)SA6,TCF=RXEZ)/OD,[T/JU0ad^_W2#.JMY;
// K45fQ^([Bg))LJZ-[P]((5K^TT3WA39#Q)Xa?(DRa&#VEGM[_dBIY]LdbBH:]1[#
// DC1>/GR&TM][)^A:.V[E]PXeP0gHb32U><:6>]AY]Z4&N;.eK]daR>M&Q&9/]MN:
// fFgSEOH=8^07.P]GC=0AD92BJY2VV-9YaL&7.5DCbREf,<GD<@_c?7TBC\;YANG#
// ;&\P@)Y[ceE;C)@??f1c;d^74CZ;5,Cd3_VI/;A##X]NKfbZ##P&6D5U=(9bC)=+
// 3:<--^/ISAJDX9.CCG9)b7I=&g.F4#5aR.K.,TOKGHT^&M9R9MLI^@AV0&@5Ea^.
// ^#N2YI2cWW:D./33LB\a/#0_A,B.K)D;2&D;[.5:1AC/bRDX/Y29,/IWd(J/a.;S
// UA46?^5X@3)d3Z\=V3HHV>_YFNCAIKZ<W5gW]>#aMZV;@QQ>VgZRXZ>D(L27A-(J
// &?V-5M<VK.Q2CX?ROHCIe>/aS:G-7O[c@A8SRN\LLPKJe_96DDR<J6^=[VJ=@PZ8
// ?H10?Mg559;^X)\>CB?8Va2RPJ]B,A[OBHE2c5Q:Y9IN7>?T\Y[U+[e5Bg\&S6MS
// /00J62gUU(?&GXZ2>Ec7-F(JWe&J)7U@=)T,2\f=1K.+,#?cHMO35F9;b85X?Q@)
// ?H[aDJB9#ZCCHYX?8?5_ML-D+EGTc/(Jf0aP9LNZ)JGDV405+Y@GbbQ.GLHbJ58O
// @5CN[D8[QDMINUfbd?OC[\#\K_XLe5O^6:MKg.JOK=#e@A=U+]g3^DFE(Q1^-eS^
// SXeU2,4G,4C[.;071/@M^83.3U[^Q3KZ,2&a<1[,?/U-bO?)]B16[(32BV:_8Y-_
// d4aOWPML@<EMZ[,UOe.(e.XWFAPQ/=H2(_fN-I_#Q#V.TZ;GS@2,B,O[6I.E6/g@
// Y>HO@\ZP>VV/PT<]EFQXaQgTEB+KW._LCfO(&QC3T7d&7R&@(TE:Wb3LUPYI_:PG
// G\@NX.6::ESGL]->UNfTL8eg^9.a6Q3V4MB6=-TJ8A,EKY(R#3afc[;3gM&F]3[Q
// :3fAGa(N@>2#,)/E5&NZ@X[VH)Y;.<Fe/\;c_R,4:Tf1cHDS#A4fba=H2]3Zg9?J
// Z:c\GU[^c@+M@]0W7cgK]Q-2X8#X+2(&)L\Kb,^FQ,:9-eT?0>XJ,K@BL=+.Y=[H
// MTT.:W>1UJNA+c55I#YN9^3J8=VW0RJDcI<6DH),02JR-/JU[&CfO,JQ&g^2+/EL
// Q3=#-@E)Y]]TO>?UB;.Mc^Z&TcYWO@5ZfQaE_6.)a/8:ZP,N^)ZSA7BDLM+?fX.5
// BdLJ#L&bKSO(\JA\A?P,?/94b2VR0T/1(Uf/WMFdK04/_8YdU=XNN-ZETaHG@U8I
// XJZC1/4AH6.+B@8P]?LCPLR2dd9,(FNb1FM04L.GPE.6K;S.RcS/:YZ94dOEQ]BG
// &C_LUOKIF]K7V+6\K_X_EBTIfFYaK.GbJ0Cc.A>Mc<=P66d<#)_8QG#VZf[eA/97
// T&C+_-U2S\_L&I?/.;?N5.6Ma_N(EPgTWCR-W\\VPI?>U#XKM,Q]f7@XPKWa[V9(
// a+RHKYF344QMLf\[FU0\4^[TI>b7<9a-5=b-M?.OZJX0ZPdQc#\&FTf&/KW(N;b2
// MDfeEMK5Y;gN&5RLF)\ZUIJO&=S6301;cHM^Vc?\(=(R-9LYMA?eaAQ,Q0-UJ2=Z
// X366:<2AgP^Z7=F5CF#Y6-McUFY2G5\OQ:)Pg_.Q@R.V=c_A26-gSXIg1SMgJGQ2
// GC#^eaT.=U9=(&#B+gQ,+f^A^&T),/[cXQ(_PaOHC&PbZ8B+4GW@gF4<Bg._&J>2
// geXc7JVVQ29#Q8Dc9\SW[#9.Q,dY)T@a25?f0KJ<A4I(<bM0IO88=;,bQMOfZ#OU
// gGAK;&d\Lb,D#5ELc;\f^7a38@ZP^ID/V,-,_5]7Igc5cUWM0L[WeHY+_Kb#7NM(
// &>E0].(R?c5KU-HUIB6+-d9>Z?^\Q2JgR,:_a#@A6cR;=bVFZLDP;8?0-d7X[=6A
// 3V#Bd&,fWU3CL)\<)6+c1/GL.H078BM./LJ7H-6YL6ZO&g@aCf/>7c^HQW@?,XdR
// OKIPVRY^=6fT:M(EZ?^DBW?5[[7Q&^Da@Bb-<<;B9fX#22.1BWfb8-(&dTGDQAOP
// S^dTg7Q00B/5I4R.BZ<->7cbO+JXJa>1@CJL,b3WP=5K\#=bHV-WQ@HWg?5e=-1/
// 7gH3F-?9fWC4U9OJF)0)+XZ@b,0dGIY:aKgF1,C]fLXI.]4T;?#@(eY#3ZBc_&\P
// \H51TUgO(EaS\gH)DR^aK8LLgSC2J_[+[]UK;DNcJabD^7W6I?.N&O[MXC(QUL@N
// ER4;_3g^Df^Q-[,bKTMf3Tf8)U,?KJdG,Ue_20@XE]2MVI#[U#)/cDg)DONB,D4]
// ;<JTVWU<O05\AZ5PG^Ndf3WP[T:-)UR.H6LdHXgB\)&ZD1CK5,CaQFXTV1YZNU#O
// a/9:#J0?c^AcRdQEdCg7a8/_GC@B@f7/bGF\X]Y<<-WR#C=dF#c\;F3<LK^Se2I?
// .?d80P;C\AL=/(;8CeYC-C\2=A99TI>B@PDg=E6.DX&a+VC:a^K2T=+R:O9-L-1/
// TYU\d[6XM-)]GMQJ.#K-;:42GCW5&[5?:(;,_M@GaQ#[g.ggP0a#7_a0PX9cc0>I
// =+#5+_LHD#@4&/9#?V7M]-D,;H;-4<e83[0.]46GC40+?fZR=BWXL#PK?HG(2A)5
// ).9D7[9;,M\HA2^CE\PWb_Q/b&b8Y6RLZ#UJ=Sg4QM]UCEc6TaXZ.ggc)2EE/\2b
// cZOXQ1d2(&2XDDBK&7>0+&FI7N@>YdfXD_W?;Yc#]@LT92P-f<(I9ORI.GOe&afd
// KQd62;+dQA)J.K4/Z<FUD#UeW_EH67>\d>.T:)0O06@@gfA>QFH_W1E:[#3PYB7X
// KEXf>JCT.67;dYY\LMb(&I\WJ]VPNWdUN3K)4JD(RT7ZUb7O&69_a5&DY:B]?8()
// ]S2Z+C7;:f?^@/bNG6WO1L3UM]+]B?fWW,1G_:6d(J8<IM&B#DL;40d<AZ8XcMQ@
// cLW;E93_]665\.7#8U:3=?8Y)E2Gf,SCcdIA#eE]>>efFX1CND+DR(5d/3C#\;32
// +1^=_91)7Q?R)gZBH&\IA:XMJg6@e>&DR@<_dB/L6:<SNg]<)3a\9d8c/a.aW@0W
// eQBCR^+QXQdb.H#L<^<C/J;>d.NJ&B<4Y^a)22&)=g6?RO9Zc.8dI:8[[D>9DAVR
// 8&U4XAEA5,cCVJ#PH]SHHV9b5X)K3.JD4[.0G0bL^9e+;4f25UWP-K#HP]I63SfZ
// /b?>2/J[PPI^c>8#R=C<&PeZ9(AC.1E\6>D8U4P&eZB#dLVDGaCSMBE#IbWcg8gP
// WDK8fb43WD>Ta0,Ja1c8)D7=[8Ea[T#LK/,[6X\D[&SZ9fBD-JS@_Z5@0Y#;LI<6
// N3/:=?;,.5#B1?DTbegYD,?Q=[YNGI6PQ.Z<Z=Q@ROdcJfBV9N.6:#aI)RR)8C[,
// 99,+_SLg:O-Z^//e_6dT6O&HgHU:GgDJ_\J@7]/LI=CLP:b4&EW,^O^G/(#]08B>
// @?d[].(./b1#(S5V?ISR^K>Ng>]f[b^1.6_4Z<2:eUVg)0CK_+X]dD.1Y?Q<)JB+
// D,TW>96)>G.\(M@#NR>Y-87T6I.C<DGD++D19>S50.5J//F(VSZYe_T[J0K5^Xf\
// ILf(<F.378@NXgFT[)g01BAG:J<Jc+\99C9)]fGX;QVQ^4JFfZJXLL6JH\8eZCQ;
// >K#2\TCO,PGCg?5aA:._^K95H\VdCYUG3ZdGD?MFUL0T\H4),])8=J0PJ3ReA][C
// JcXBA7ZU8NHCH:EXF[8M]/6XR7/[?[A19X1J6/35LS9&[1Y]4H1P@-c9J365ZBa>
// <]N6:M^VS/K(,1@;3TdfeXbfG(^#(4P/^dc4M^[:21P5D(I,_b6Q@>-c[>6W5O[N
// H^L<D_B:a/CAV&44^PJ@d:.2F;fMCGJ8DAKYV=8Z;d5=#S\+C-Y9X:DRO(2f(Lf8
// ^#5N?I82=+056B23GWdTFUbIaA[FNg]:E#UOY=ZAP?@BeG:#2eSc@[0QeL=Sg4eP
// Z85f;/1/)+?^H9AN.+S)8[JAD163<KYMNL@.62YYX<0_A4_<1cN>Ld1,A1WEY:XH
// _d=P46(XG6B5:3?[R91^Q]gcc=331N,;.]:-@T?S/A<(H#NWQAUA_L+MDOJC_OCT
// 9?QD:ZF::P5C6FC<(?2A+(K[Y16<]a^gZ)ef/AR+1)A&<^&1MQ\)CEVA.I&fH(YY
// DYC1K;gcOE?6F;,Dab&>WYPP,8<8R5-I?3fgJ7T)#>XV0F<:cW5C5U>#RY\1fW=S
// K?_XMde=MY0.1+_UWUOXH5456dgaQ..7@J9g\+fD3Y^+0,(OCgPBdP+=f5(QWW1<
// Sd:P@;;.U.]SDRVBc2C=Y+EF88L3D6ggd;Y7F^O<4Oa&@>9Y]C[<R&55:d/>dP@E
// G>]>XSZ_P>5C\&N0TSGU)PUcPU(4?7C^:FKOHZD9;;EbPfdU7>RPAH.WdVH\ZBPK
// 2W6509A>(Z:PA>M=U[,4P?)&8QLH;I973\0(E^)#A,RYZAbe/H5&;45V#Gf^G<2f
// X4C>^:d]/6A(a5Ge?cP4]Lc]H<.b+JbINc:[6.Q8CRI<LIXRF:]OE&YMYN.ACT#H
// a.2;RN+7dLedX3XPC9ZLWP,@7O>=_/T9#IJ[,.D,f),1:)10[J_1.(3]3O[P@Y@.
// Z4W/DJ0>)RJ/_SKLTH4>RKHD.^bbE+1>TQ/NdR?8gA-KDe/(HJ4cK_W<Ie8:LdN9
// HH7(DOd<Q_b+XSJW4O=\NS9#[EDLSE2Pb51R3=:cR33U9<R^E,9:?9,LHCQDD1M9
// >M1K;P9\7)2+:VA?79?Vc+bgSLM\5[Ee.2.1cdbLC&,<R^4&:;0#4=C7]&.^T9D8
// ]Yc95RB7c1O:B;@PGZP=?M9-76D<ZA_:@GgdQe\d=JZKWKWI?F).#E1^C5N86f+a
// C8c@EROPV,Pb^P-1Sa6?@PbdX,SO4\ZSCedO-@-(KC-9Y^J]0dBE4X@Vc+-C;/g@
// (dRJ4^71;AY505:b[c>K4^NWCB/T^:-SET.G_U>:(Kg,NW3@O)T[IJJ?..43U\9K
// :R&:Sf(:g85DdN0JGR65UgS3?QXG8>0B[U=9]\C(C+I?-;XQaVLDf@b)e=5Q]AO8
// ;-E5TV(5B-N9eG]Y:C\K?[RQ-W,c,1Rg==,dG6IPI82]\d,+,/+,R<?#Z61aEaO,
// _&_0B1&0b_U<21)[6(4J6BA@J#eVM.(aYbND/[5FVY6?R;C>;PMB?(UZ0,S_I,8T
// <D.^eI2\d<eGO,V8R#:ag6H3L8-RTE_Z->YB:(7.c][A=_c:-:Q8&DVWP21g[)f^
// NdLI]D8a1f>-3+b<8#Y7R:9C(-c2fKNB.FQ#&Qd@b:,-^W/W=Y_?R9WbGLfWC;O<
// >\KgT/QSM+d>F1_g#.33?^=b>0]>=Lb+BVY84KD,/[IC9>)3=R??g,X2cbR(#=E4
// Af@e:J?+[eZbJAO8dV>e<<L?e1.>@3#?9RYH1NRgRU\#\MQ7eT8#ED0(,7;[Y(g@
// ^7ZI&b,f&HeBOgQVJ#R]JOf2X24#J&IHC=f+SfWAB?7dDXN4PWI4B/>b[1(7_.R.
// N8/TUD@(Y@Y+>MLBD&@[C@R&BX)U@/@+e\e.Jfg>VW@af93Ufd,6R2P8?CBO_]8Z
// )8JQA6=TZ(JeaR-V6#);a7DRMPcLJW(.TD/6^8R-,e)cH?F@H5U(P^(6K6UCGOZc
// WdBdZ7^I&:Y_XAQf-cYS4MP3ZG2LX.?Y<-,W(4/gVPIAWJQ^.COYT/,<F(72BEKX
// 6d_^I\S;eYZM>K[T76P]+/2QNV1WQ5/4Z+b-596K4_L\[A[-QNM&ZW#ZK76be3UQ
// JS2S0@c,3W_O6A]12LAB==fgSMT>LaF:dALVZgNM#/9+9)AV3AFEa1W^&QD8]MFN
// ?@TG.P:K0Aa=@TXC7=NC4UO:ZUcd8@#e8,AFX-OTX^TgAT<QE<?cGN\F)=?^76ZY
// R.(K_;9[V7NF)TAgMX=H7UE88-a@<K44YZ]eA4:T(BN&23U0.8Q-Y+3@X3,UCEX=
// NP@(5=DJbSdV>C8Be7+N<:P.3f+QE?JaISQ;PdTK\5@;L,8FY(fLV3fAGRBCKVE[
// a@(c#/;KG784>DEN&d16AOLbd+e;T1/5bcK(c0.#8WgNDL0.ON0>_4c&fW3T/#(Y
// J\]gWX?2=G:Cfc^)Eb<=ONB.6IB=#SZ.TH(@aNBd@WeOOHgXXOTE4cZTeLPMNgTg
// :C/;gaZc&PJ_<d0N31gc#JgCgFNC/7L_NG:>2^-af@(4-LfT>JH#B6PSd;CQ+^^W
// U._I==J28FFQdde4PH1Y[9fJbN6?]W1<0J8?fgNc:)G#HEM7^Cfc]fP]OSY56e8g
// ^Y0H\>TgB\W30>\6f)bLL7PKgf=H&P<523XY]JcGJad,J)B>=9X8.JHN9?)Y#H7-
// 8RN._/GW0I>NgWP>=^D?GXVPBGXgKISN8O[3VHGMLe+9>43,H3NY5S0WbX\>#Ee\
// Q>4OPC6b68?:M4R>0Y65_SJ3E\cA37gL70CY]XcK[9)+_3B2AaQ,48],IDSOc)=/
// =R+ZAHWbY[\@6)GM\NH;MbQ[Q(g5TLF9EA^8g6L8^0c\X<(@CG/HHW>@d+V1@W5=
// -W:\HW_ceaX\_3G/J5MgD6BaUb1,((dRBVKP9=cG5R7M:d0^M/+\aH?bIB:)X\=Y
// M;H5TKW8fDO54FZ5O?W.9@T:RTdbM(cIJA7HEcEWWC^I8/HaXPfaJSeWb#fQ:e6>
// Kb0@F>DH)XX@7=Zeg+I5BFeU:-W<6d,eZI^Z-a7=&66C0P^D<LbVC;#-=(EgKZQ]
// 80.N]fHSI?2NFH#e56b^/B2;VVfX)R:JdgP9Q&0^S1DZgM.-,[a=VQD=)8W?D(de
// 1]EaO5J>_VCXcCTY<K,I75Y]_2RVE1g;eYedE?(/b@X,.4BPNK7a0D,J,WZO4gaN
// ?\eLTbM9][S2<b@FSLg;=#A+W,eC0-UeJb4MVNSC+>E<=/^S/#H=MZ_:H0_LAf6X
// 7,L,:/f]<C5:dFJfU39;K5B.)./SCCI4#FD:;ZP/+R\9-a]IE9&#.P/EXOBET\@>
// QZ=7S.HE#dZdZ9Y,^0-P)Y[(#]53B-E3?O?:F;)LBCYB\DU???gYQ^?8M?6);K(&
// I=^&a/(g\U)>-2aOPXH)-);A6)J=[Pa#+=,PF+U.K_He\.BY(FMa+TH;UG50I5Y<
// \67O:_NQBg]Q9TL5Hb]c]5d9;R1Igb#QS-)LBUE:41E9.<B?OBDL3CMLaP,,@@MW
// =4e\DA:9aT_df:KPM8+Lg;8NU^aRXO[#&F22GC^bQ>&6\2K?Y?&R8&08=RVB\:6]
// gU95:d=U4I2HgK\cAN#Y)Q_85<:N4KVYYCIRg3C:Z=MYUR32=&KQ(fT@?GEI&C#g
// >+OPUXX#)\PAPS,b3+[36LWGWJ?V&cJ/>S-@6/2S6HO3;/?5@94[g\W#?R=Hd]J#
// [EZ?R?\U=BUdI3<]&]ZQ_24[_BORA))D;ZeVa]<.:M>+BVJ>J?c?=BE40)QQ:UQ9
// gbSgX=6>4a+77==[;P2DN2BM:@T/1M_::P0f6ID9TV[-OI;69BK]OBI5gUM9g5+A
// ,QM[?]FORT\bN1E_]M5Ue2U,]WBBTH,4M\cgcX5BfVHMgYX9PQP;V#IPID/9MZ]F
// L[N@AEE=?[NcP)f^:W6dg8c1gUEBg5a6BG1E3/?4OEAc_/U:C)(LNA4G-VKNY>-J
// 8GR_?;8_>M]G6a/8)V8YLK?N]VG+YfYObTCCT6]0F75NWS?(>S\DAcLE[F&-[e5d
// )L^:2Mb6)f6/LN)MM[:5GG]EXM:HbI3L(HD&]\IG9A=JV-^GL-g[Yad&]P=.^3<4
// FSg_U,e+^bbX:CbaP2E6M;FO8IZGS6?^Y:QdW9.aS0fIg=39AO23UHUO,/-B^Y+/
// 7,K[+RSJ^[5Tfd@A<O<P^-MW@B_cI=<aQPCA9TI=H46ge?8c0:#[AM:])->fU(,g
// >O[gAUBPPWLe(H@SM+]20.39:,2:5/YJb,HfZ4BbE,]fIKfJ@+5^/?8.YL#Y<U-H
// JIQ=,>;98=;<IH[PJ&6<[\(WfMT5gI0GCdR^B;GS=ND?9>dWE3#=;b&T5b>7I/.=
// #1-MLKG/bQQ#<1=>?3WTO>/N8\FdAGX4/[THXILSO(W(:+L:I@7A)MQL<>TDVS.a
// Daf8]UY_\2LT?Y54a=g4)G/H.E>:ZD&6gAf.g/1gJ1W7<JIRV<\>3<(8_GLN768e
// TI[B-K9RCEKN48>=VAePM5Q>A@C_P@gUJ/>T6Z0V<;OJ[CJ:Ae+WdfT;16X,V^>3
// .(;V.eF)#Ja<8Z9PgE9O@+JdT<7b\KH-L>T?6,<d_GM1249fO9TFJ<>9)#?X#FJL
// J9R+P27+X1?2\Hc).Eg;HfEd=E>a@)>(TFIX1U0G:FW&A5YM4eT_@]5]DJ7NVDOM
// 9+<WN0ZN&IDQTd;#f1Xg[WE_>IFb:J@#fe2TF\WD5ONg;?75V70/K-]ML7XI]0E)
// L3+MTDICK_UK12&2J#(=2)/M&BeKg<JJYDJ<Rda\:\1Y36.P;@_6B<@+ZFR4Z[4G
// 8)2f;[\5_J1;V(A9>I17dZ@10-3]0C[BOH.,PFJNAARfVd=CGV<3ARf39&4+@>Zb
// S2@UPGSHD404Y\2OW=9eZCU/JGK3(-IV_M7NA-WF7P#?&9]8L(2^^H,Q;L>bC^IB
// [)eeS@\/-FA(B[2ZG##>Z8X;eeOG9]?AN2NK(]2Zc95Z?8+AD;+I4X15/cN7MRI.
// I_>ED/fedELYKa)X-FJ9HHD/=LE2G+.<gWU0<PR=O_-^e/gU__7aJg4a7Wb=d&SV
// L,/3)[5I1Hb,ET0cOJTa>?4)86bY_6,ZN/9#>?W13G.34\;Qee@GSY9LPfMR2H?:
// (Fe2RM6Rb4M]fKbLW];3HZQfUGBP@b,>+,\52<V.JRH-YfMWL7f[RHYX1ae()gLV
// M0JbQ?R1R<WM@Z+cTZRN^XEU_]\GT_[RVG@QFHYTQeQ-bUKWUC6eSdNMR)H]1\;C
// EPYgCLER926]9V+:a/DUJXU\.D?F31L0^@A.)\bd2A>g.-<T3)0UJ3MG;8R#/DIf
// b/Ygc<P.-4H:&7Ae5fW4?UISB1<fY/UMK8BWNQJPN57P->UHEYd^8F_\+7EZ2.62
// a8/R5RDB+A_&WY(P>e66Q]FA/Pc[W]>3/1^052-JWId6S,V7V>1;P-]R8RCQ#J=f
// SLJ_9gV/3I@SPQfbN#<K_IEGOY]Tc(W13]W^^g5WN)A\\U3/I^<:M?NM>g.AXc3[
// N1a=0\J0/^L&E1C45[656M=I;#4RTgdW:9bDWb507=fD_bP)Z8(eE?Bc1c=I]#RB
// daCD^AQKSNB3>;[N\DDcfV48AGX1a_S3Y)-.=N/DG_5:d0Y]Ce2V-79->K5DF]fC
// ;BYaHK]d[S?+8Ue+T,E\28#7#MeJc+QH9BJ-=M:Z.JA3^IY75^0fg[EZ44L;e^R4
// 4D.(WfSXSgUT/)6<4/\O.&:1)OO;-UB&_=PegC:IRB[06F\YSIL#gVYZJWE]W^@4
// \ZPfdg]IU.I5\[R-,TBK7,cfITC[N_1C&LLD<BCg6b<73L/.\E9J@=:9ER#7S+_P
// RO9N8]>;B>;eLA#P;cX\H<IZK1T:OKT##CO-^E\]d.U(TV6F(P]EXd_-J6J;>#[_
// #FJK(VE[)3VWIS/Y0IQH/LXKA3DEIeC43<+;H#BGJNZ)1+_>A[3TM+W-GB#KN;2P
// 1(cS:9?7bQU(?T\;4d<(>_4V;0R7HAD9g=Ed\A7gWCScWYT2=K30&J5S.cX&,>3c
// ^)_gSLGJf70+<1b?QG<,[I\,(O,E-gN+_;LW/539QI^BPYO^Z@c6]/8#8a:]Z@8#
// +f)VGWX@1^),^BQb[JeV#eIC#I?0Pg;e]@SX8E,QQ3c#fL_bLNcJ)F5f9R9X-U4X
// 4e7F^-2HUg,:G)^Hc#fVDb3b8RTCVb9,.Q1N<DFgCQTcdf>^ADEW80SD8683eTB8
// =Y<,,_SeG..2I9g9Vd5,;==e[,gFgTBcER9NCKF\0LebWAVCTNV54DU16b+OA8@K
// 46?aO]@-H9&Jd.ab?R8e2]HJd)U#FJ:E2HG#X4ZUa=#U)>e?3_<\9K[@JeQ:JC=e
// )#&;#9-#G>bEE(272H,SWN1,08^(_+K&R;=52e_@(]8-W?#fP&edTbAc3VU_^9VN
// GeO6HcE?@94R,5J[6W2(PJ:]VCE+<dY4H]S=BXG.;>0WHOgG3Y.Vc#Pe7839SA\e
// A&YOWSC-RNY3?]=5+BY/[FW^-gd5-_5JX2(P_S=WK8V:]6eLE>=LHeb>-P3.2_L2
// RV:M-,E8f2#f8Y>RNa2FT>B1cB40VY7PPZ+S90CV/>dT=Fd->UQY&[-?8O0gI+KR
// b(22)/F>A>)NG?6^b(4@&+5GNX.gX5U(6V4[E&-?7GWWT.T&>K#A3-;363:04^ZM
// g8\eKYecG[5?(aNZfX::Y-7-:KGg;;^8D>O-9]PHE-DLc](IX@[U,YBG&OW.IZL+
// XNXP@SJSNb;#^)92@3(ANbLD7JQaAB^:QHX@LdD_.cXV(F;J9\#3.g=)HM[Jb7M?
// FDV<(AVRd@HM@OUZ;TF[&6_TK/\-M&LIGaLKaOUc^S2&=<e2ebKP(JXQM@9SZ,GU
// -X)G#cE_EF^b@3@)G?)+U+.IbH3Egf8?dGecY,:UIY.SIWDg\WNBR:PKH(-CE/,:
// K)J)0&98>C[0]O=7UQ\-8A:L+QVbbY2a7=,eZ.ecf<LV<dUE5Z)GH)P+ObC_?-60
// D7FPCg?0>_FVg=X#P+f0;V>7V/BNM63;ag4BH+FQ[4K\Y>N\dH9PWTC@NIU#1<T;
// G0XeG#bB=R_/)D-E1Y+>E.TAY4gfa84C&:W^1<8)9HID-b/1O.HVG=g8(?V^BH-9
// PEB4dNIa^F[a699]F9FJ2-0,D+_]?E@(J2I?Vd1B:_7AdeRNWD;J3?g_</Ue#J&:
// 6GWD=&_=>d>DL])TD.9E]3L7T5;<TU&f[#WT35RLfcXHU.2Oc5F^Q]2CU?4#+2.@
// )ZDI@JK:/+WK5.TJ4N8+QBWG4b>[W:Q&ZXM)-Xg@/?baYg7<<^APE3B^##>G.OaG
// aGL5CRYUG9T-9?E6b^D.X<8CV(KASg;]Q1LBJ49ef4K65)f2+:#=T\;45a8^N]K]
// )[ML8L/B]^ZM&HOJVJ/:)G5e^]8.64+PX^,:2-&b=Q;\MXCVAcfK1D[4P(@S[A&V
// 2-c(:ffBY0[,eN2HU0FRe^b:,3B99(,Md/0@T^/NF5V8S)5f=Lg89IPETYNc)g4D
// )0UMX[LPNaOLYa-,#E6>/]K,X(#DIAWU#);-7e-<gaT,<=1UQb@+]bKBHNdCC?_]
// E4AP]3)=ST.g8JKRI]\.bRW-PE9L83:QVX0KIK9[cV>gdV&\cQU,E+W7#_D:2#V0
// >=(SWS3RM79VB[8_]IgO[25@fc12KXJ=c8L@fU0TRb3&20KW-e8)Y_d_&26?P,W]
// RTFZ6BFQX>E?;)bA]^/>9TQX+/X;Ab5.0E,VL09?5,AX@<_G3V;cOb?7_eR,2T>G
// f<R_KYBX;+V>NKMB?I=Veb66Va,dQ&>\,:_YIWcFN:c#f[H^OZS]c\H=ee[_:NN#
// \LL(X_4Reg^LZdd@C@a\-CCXZ8PD-L(^F&N(R61:[FaSH]5FJgN>c@U0E0^CaeD<
// )=]^(T&=T?,&_8#O;(Z8LM/2YM>^+_:XYKAE;?,6a_GVbF/UD=J/d[(H]TQV\2;H
// \W-?5AB:A)45a(YOT,@CE#L.L5[^6dG0c7b[&TRI5,H-/a@J7FPYOdG6FWZ>R\]G
// Mf?+CPIG#Cg+>:F;A-C\g8[eD2QX0QY-J6CcWJf;7Jc]AP<1M5X16[IAC8I:B+@c
// cN->M_1gI#_>VXed?)a2bHMF&]2BIH@ED7g1;3fB73@^S33aV5@W1c)MNX.)(TY)
// )-[YV6K[A3O0).2E#)>JNeOLLJITd#XX_[AP,>f5.eIU+B7[K6fMf84g?I<#+5MM
// M-Q]W2XT_?@^C.c;^8_,.IgaQ0U.2^e,^2XX]3V+3-,@bAH7N/d6==^9.?42FdIH
// BP.<,&fd#PSGF)TOJf36_@B&g;M_=<K6WU53a<L:E-I>Xf<9Xd31T5b_3dIHH>I,
// .7?B8F/Q54EbEa5DMQJ?^d11G=06W=O6V/.H(WHaI8aK\f^4Q,YJ(6<7OR94UVRP
// WQA&HYWGRcD#9d5=B?T_0(e5LJ(#HR9HK#U\,=:7?H6;/PSAYO\LYC/:DWc21a9K
// +4(&CZ,#,IU>Q2g9-S-JRXMEQSW^6ebEI+M_a40.=08+FC)>d(E+3>f@U\T.7Vge
// =68_/^A/2c0<DTdNf[5790)#MMgf]@/]D0PI#Q[./>E,Ncc8J@)[XH>V[K(U[.[C
// EP15II(IZ[aLFfgK\^T)&L\1I_)RQQ#H=c3V4.W/CU@;Y2T[];<^7ARCNB<K@/8g
// gWR/N;(3565SeP.[V[6F#NHP0G@EAc_K#/-:B,QDTA9;_E[:]F>C[P0X<a4C#GTX
// \1M#1g17<6TM\82..F?;-R@J;3WC1I3UUOCZg>aI_>:TNf[AU4XSb:?P;=Z+b\BP
// T=U.^6&M24TA,>1@[^3ET+\cP9TbT747)G3.DW5Q_R,,eE2W9I)UWeT#&fWaX&OI
// 1;_Y,)dAIB;-28^0dI\IWDB1]21fR,>Z.UF<aDRAH.?C#OC\C?](#/&L7-Wa)a0/
// 2eCJY<Od7H@@5@?2;\&+(SZfZB6JSeJb4bGJZ(I_#[1XVI6c76f:a4NN3bgX?V,?
// )PIH5/GX0\ZGRDJRf@:4>E0[U-c+@6O1?)Hf2R,#c96<A6Q>K&cJ&.Yb:JA0b6/5
// )0+]<97Q,Ab;_=UL<gEgIER<DZ6@:1J>4L(D=f[NZG]9e8Q\>UeSN6?fC]VRXNL5
// 8[e7^V=Z:C#:_QQ8#:5P=KN5@\g.LMW5+,@IOI:Q]Y5MS<P?@5@B>9b@?EE7EAaY
// [eMV2b@+,VGg57(UDOT3Y6YM]X@d+82]YP+bFYfMDM+M&_AQ\KQ2:(DAgGS#PJ+2
// 0U/STMU9Q[[:0WZ[SgMNZ8a>5@6@_JK#I\a8GFb,2F0IAH9_;&B<V]U9UaPGLCUC
// JW8PG=;b/cOA2DJZ-dI/1=AZ^AK@QRNJ^1K?1L[Z[\FSAWCZ:b;+A(,_JWQLRGLW
// \ZUbe(c-5/B/NNW=KBP)DM1BMB(NE3MN@ccS>^JCHJ6A@[8+?T=e),M(G^7f:E#4
// #OdO<3I)#bdcP_Ia-LGX2<3.I:0H.50\47Z@Kb8ffdID\9_1P6Y1>dM5G&bIOce[
// +cW5K9I1PH65cbMe=)@[H5Lb?eL^5I[HOO4)A]M0AJTfE)@(;CB:]g)>R>/<OLZe
// DK]@3U75/I]:cQ#JKPV1K-2SX7NB(Cc+1I/Y-7C27F+_0M(,W\T(V,@+P?5<C)&c
// bP=+@>A+^9F4dQYL;X2@J#F-)/cCO?EFfeZ-5ZQN<2F0CE74e7cK(#A(0)88^JMP
// E28F1b\f8b>X#^__154bRa:AAW1O[M/,YFXDPEXQf1eD/2J03[N--(.C#>NLfWG]
// 5TebU]&=<^-Y7IOZY=g,ML10_O64PEfF8.BE5cbS#J-2>bS_;T)J]:/d[IVf[_<0
// ACPZ<36E8^8L]?\ZE2=1b\^F:-598;BgC1a15&8fa>K#2&5:RQ7TL^LfEEX@A,C(
// 8>\[1Xbd7FL3KFaVUZEAaHJ]F>4B0QBQ.a?Oa<LP^U)F0CMU#5M&<ZKKPS;1ZJE5
// WC#RK0Y2(g9#D^3H.>F9[BTI8=dAA(G9?EDB></f36#=<:P)\#/PQ0H#^3[#0\US
// P4W6SI;@3E43Z@5G)(H>\[8\N]/ZTAX;QAS[<_NgdMa2d^2#3/+<Z]?&>?aRMJ/=
// LfeKS,DF&L1>;W0?DfKN,Y&BGPKID\10VgZUVL0I(H[<a:.8R93#[UP,aEZ-b=>&
// 79Ng/C<3CMQd->ccI;Z.E6(+@Y95WQ]R)-Sd\=&NK>X1fKJ1:MMS2E\)_-R_<&aR
// S0DV_>LSU0KQ;S_DLTO6K8N1?@QI&/cNN(Z:5f=X&SS7B@b\9N7:B,KZ(7B\0HT=
// #+A0;XVS;6YI:Ef+3E<S&g]c)/^_V2J.:[9CID@#D7>MQR#CX-QHAb7[019AdWa-
// J^AdN8bdL-8B]73CL\KU8=gb0[dObDK]L+2>GE54V=]^Nd,1]V5X#+W,>>OBN3?A
// ;0]AMLG>aVEI8RbKf4Ib&/;TRaP(Ue]6_[d)9NUMD2O1^P16Sa609[-;2e?Q6-4<
// 9^;U3E=JW](&AT&X.;S1bWM1Cb:S>a:@QY97T?RFS5Q/ZXHWT+J>?HOADKTL,H](
// 2H,VT@,C5g9F371XQ,5>/OD>Ra#42=AE)R9A</7AA8dYFISC,N/Q:<3g(;M@:bb1
// I)(2J8e#<(UJca];6f:N]Od^d8?I>KVf[/7_R#DMJ4@5f?HK]7;ZNEA;:6U.6S;P
// \Q^S<:_P@f]@F_:g=NNJd;HfM\MB.M7VeaS8OOVE>VZX(G;MUdYb82;1@W>)75(C
// ba]:Og0^ONPcMZ)a-A&.4)\.b0_>\)a=NMBKJc<C;)/IG6-gRMBe]BbQ#Q13F6BS
// [3OU);M1.[19#V45;Wa?I<E3452#7M\b+_]g=7+W&L\f2=+Y#W81dIC[7bQS7)9[
// /1Q.4GQJ-P>b>9L/&VC+U/=RJdTG@(&7+_C>+4O(RZHUV(GDZ@ALJ1&G[KR+AGBR
// cHO;gD+Tg=G1&b2\GJcW1ZF@c@4c[9B>JIL(g4c,G:N_.TL_E^.L51D0DB(@PG@U
// aOVE38FE=bX5V(\K8cB2=8R<;5O8C)]Y+>K0(80NgX2X7.1H-TX5QRgg^?WaD4-W
// H->/CSANb#41>:1e.HF9c?M77@OGR56S(3R7YE?RTU=TG?a,cWbS^I5/ZCe9<c]#
// FT-/RYK.Ka9>DW/&.(-);ZCR=7fD&cI2(_C-ac?WX:?QKa/N&S:LCJ6D059J&b)F
// VKd7V]fVfYQT1K2Xa7S\1HVC?_^6AeI)-1+g\.&2gV=2=FDE^\E4L5-3JZaBY&3K
// >;+(M@VM=4_]2#EIR<Z2SeIZb8T@MH3.BN>]X&JYVLQT_T8MBWBb/;MTSN-3,U=#
// +NLM-dI#0Y_b(AeJG2NC^9OH()ERM8]RZ[^.Gb28T(EV#7cOW0&IUDZ=[)X=6M4E
// 10NV@;5aK)4<4(P/X;;=(=9?\+X2DD_G0CL2/&JVOC/Y[7]?5?_dc,D0NJ160JQe
// f(R52.a<Z>=DP&bE6?Z<S8Md,R.aM-6f)<T)RdVf,7,,dOZZ#+)X]=?K_.J/\),:
// :BM58>56&49WS[J[R<ga29729(5]Q=Z\e.,9:b&:P=I2+V4cHC.XS34<FCRRN-L(
// U=^&[Jce\\#6R>/__&1D2\/2[F\eG2^cb=-PgK7OfLT5#Vbe-@K?c^E\8+f>XCDf
// BXOIY)e^)M-79>fP;+N(d5]?FZH[L]Z<K_Q0>>AD8^74X&_TBd1J6NfB?06-2]/2
// a]aeAT#AVZ(3251e;86NdYbPGg4D12<TL;41RN)eWNO5W7E4VHQEMXM3P;J\UeCX
// P.Z@AQ@=.9[eWaT+-),UXY9KE2D],eJ3\INT:NE/T;+J=F?4L4RDgB=H7c5fb2(4
// ,7@D,WNP0_G?VT4^JOH42B)XQ>H_K3-X+7YH,Ue2&/<XDDWV>FO18ccdA=9N82K.
// ^DC&HH@9V:Hg:b.g:7(_)L/gENJ]IJd^^Q,[:CU6&]\_f+AV1^QE-.d4X==TUO=d
// L7Jf8=/<>b26g82N^DC[32,+]>V-[WIf0/-ZI#6954gcaB,):?6F]O@LH5]E-1ZB
// KT:P9K<WUZ(X(.245SD@3eHeF5d=K#>2BdYRB26.-:&XX@-H+F&EgU,2669?\TE>
// OaQ[P/UDQ,LQW@f0?4B^C0Y.&&\F_)-8NMZ#WKb6;fW.^\Ha5>/G2Z,MC/I]T28T
// J7&fbF1L>G@W&]@5/aPG:?1L.<@5IbcMY@8Zd89[B#0>3[L7TQ1WX9]]W4J[Hc5>
// 2P96V[LL4^e,?]N;S(-J\Ec^C0[C,=-[\KPW@K[8IK)THSWR2aQ:V1+V9Z2(\K@\
// QHXJgJC]gf+MMYKS?QB4?J?U.7:/DYO+=43ZWbY=aNJR6f[\+-#_CM?T_0Ac62bG
// b65KMbBA?EeLHd6=3-PF9,#0G4P9@2.\UCU[>KENVOXYL\Fe7K;CH^Pg5^78=,FU
// ]H09#SY-a&^\.H\GDC#IS1gO1&#W0K>K,MUf6g7A)FIf)Re#+UDBHYb<QAQVC-&A
// _W19,Aaa(bHI--TI\M[&adN(1:G_T0+<E5f?7F?ACfOH:GD\Z[I0&<=K;A1N3[C:
// ^C+1#\+[d(AIO>X1P0UQKTEO,1X\Z1&JQFDb-K5G&F:>#Id7;9BBfXK:9)J^P]ND
// R+b]Kgd:03T<<-:8^:TJ1UU+ZaN4U6><Rec3a:aN7.[Rfee/WA/6)aDG[JLGMKVe
// JFYBM#V<F5JN13H=H<+Rc&@PG_M3HL(E/FYYOdeKWU6\TZ2#JgaIFFQKRb9W(7=W
// :fa]1^):b^Z;9bMd-/H^.df:.0^9]1+bN<2N)0O_D/6Fg1+V/G>+AV;Ce2C/,EG4
// :2UDPOLb&_\E)J3[\@6@6d4#<>bgf4B?-;;[6(;SR?&RXPH-@;&UEfWHYE9@JIf4
// W-5Q[0(6TQd_WeI;0&EUI5.<2Lf,d:e.@c]D7X/F+MQ4cX7/5HLf/GT5^a]MF2?>
// 7\6X-f@J+b:A:.L._=JL)_.\W.V1QD6P-:NGPE32NT/G9Q=J^&2AaJO1fbJM307g
// &&PaERD8^X91I,I>7N.O4CbUD8BVU_-6.6YK@8Y0)E0#/TLe41-1=OB.4cML<5O&
// 9933V54ABP+8f=dOH76,XDAALYe+Se1>L-I((B[7U/9R8^G8G_WW4DF9FZd+e3;]
// ?_<U>gU.=TVVJAc3UI?DB7@G_<W<<AC+TJ1RWe:AdSI2g/\D9g_Z4ddPTN-L65gS
// Xg95/[US1\cR6cI6&g0IC=_>SH5]bebVG;O52e<&d\3d1bNgLW9f]LcPY-+#JP\]
// -IZ2<ScQMf&B4FB5,^QV>ALTfKX=>).EbJI1(U:E.8X-V[U/&XXX_G1abBfb;FBd
// JAUT[^[BNg+B\;B6.)VN_S(17X+Fd?QLf=IfEJ[5Y,M6Dg=YT562&)V\dR__9\R=
// GM9/Q2QaHJg))-0-QgVGe1H4/.-;Y=O2.eXU:,<V1&@<ZbBC#Q_Q5C3R9\5>,_55
// +aUKN4g1I7B]1O<KH3Je;[Z_Y+6YgA#g;#D5G4Z<aL&1aZ27:[BS4?F6Fe9TVHa>
// &>g(e&2___]e2-S5&7+#XfgTP5#@-dA>a9EUV()]gML\RA7NS\#984/;cO]2PR=Q
// YSZSEJ3YU,Z=X7Q-=QL,DU0,M9DE^NMS67^I]3SO0N[Ng(B:(.Y#g>=XEb^T]fB[
// PKAI:O?G_?QZDZaBU391\ELIE?TM7-aE2aDS(:IbH<[e]#T&:BUCQUY_6(E_IU0.
// IJVb/P9BIP@;cd2X^EeN>NbFbZ7cFD]5O&IQJJ](ZKdY]/Y(YZSSIb2;W9T(\a?[
// LOH=_=dX6RYP6BX9_ET01/PMAW.2T6G>=)\32,=FbY6eVD5,IJ:;c?+JHX/fV4ZF
// FB<K@bKg-#.@5L0L4NbM];[[HW3AJ98CSO^I6Z_TI[7GS]RB:2(9f>]/19=H<B^N
// 06KIPSfAN9AL(=L-VdU;+HDZHP1fNG4TCYEccWcc(R4LIOLW#9gOVVKBdCKag,9<
// b+<aJA,>KZA+TV6N9DI/Xd,&d1>W=UcC#]O(=P@SaO(BJB<)g3e2Z8,Y3<)bZg22
// 7PHNY?4Se80gV+SG^+8,:RZ.)6,cXZZ,BN>8J4X>_I?N:ZIKa^TIg\XUBMD^6g]T
// Og2X@gf0:+IcR98DI;fYU-.Od2Q1UcAW0>VJd3.34.)1HRKGG42@8<9U@XBLPIT?
// gPB87_O=3TMZL(bMgG(9TKM9:+Gd:0SZK3&b?(Z(U]GJ,G_VC;@17Y-@>dc^\[#a
// 2UIKA=O?c]F-\K>>)Y^I33Q[NH/4>b-\>Lc]H5?E;9e?=3(_;Q1G_eb8-QD;ea8[
// g6BB@X3YO@&RYI??NKN1_]2[:B&<XQK3V[:^e96)L,K-cAUc<,FZP(2Zb5\EOJOF
// 45/2H^=[^1<U37/@:5=I31GfO>/9JF[YXVQ+/5G#&APg#U1#dLC:T7_X1:OTH.g2
// 8I/>;EHL3bc..dZb\#65e/LgRR9GObV&@9)@86M<A.eg6X^=_),JgGe>F_-Y:#bA
// F3?cAgMD]g?GL0/ZfL\M#9Q#,a##LE&+FHYVA;_C^N0+D()2\VLa^304g:B^QHbA
// ?K3P17M7+U&=,7\BU+VDODU[R^NUEBV^U1^CDF;C?-GI&gfOKWO8Q;F/X0(dObG&
// \QW@#0Lg[@U3Y[+;:gI9&<AR71e4@VOf>Z,ITF:#a4-N^0-B]S.O=3(c4&\4:3X[
// 3@-.SdVOIVX@Ob^0(6aL\#1GOW9]TdDWJ.4.IT<&&DI[45aP]2?580^S-D[+VML6
// F@)LA3U(TPM02U&Rc;b(A3G><TE;#^6:YQ<T>F&f8,(QRT<NC;bV&I_PXR]GcG.X
// O:EacU0QAfS;aY3c0/A6_A=<3DQ9:NBAVc[g,?>B-ZD@8-fP?]KY_AI-01#RR,(A
// PHJSD34N6OXRegD2,>P?V]aXBf\R+,5#V@aJZIOc0JR[fX9U6.<_T/Q=/3cQ6IYT
// 0cHS.C4AfP\SND2R2D14U;cD0#(V3<Q</#GF\>>I8fJX6L?EH3;WLSK1<AAa.J^f
// 3/]M,7DZI_YdM+76NX9QQXaPZSaI56QB-K>@=g&Y0[ZRIV6R,@@6O/JBe.2X&IY1
// -)NIHT[>7MMZ6#4/CSRNb^?L/^UL[#>6K:@#Dc.X#b+7#L3.[2aZ[XS.6+TRD.S5
// a+JTM5QKg;(,Rf?_-;S=[Q:8_1eL4C.AC[g9ABfK;<HSL@VY4,0DGCHQ#^1E/RZ3
// 32c5[eJ)_Y7&RV4QBf7>0-,#^62VfcWD941?G]K316;Xf8#TBENTUMRMB#cFbJQ=
// V#XT[@LG5Ce1PRT+I:[IK&V=6P>POFDgC^;<J]#FPB#.f#^6]-J.Z@2=X&,I8bHS
// AOag;?(-Q2;QE(97PC(.O2F2H\I(9/V<d2VC_\a#499E#Cb9<@_9^]Yc7VC1CB>:
// R3L?M.6P2-0S0bJZHT<4dc;-e.KWOL[TOcDLGDX3AQc5&B)\Q^BI-0d06_XQS5\?
// )LfPEDJ[_Ug&+2BK9@H9R\&,g6Dc1,.61]9XM2SYU([E:WO)]P7-\VJa<>)>P,Ua
// \TbB&.SIBWWPWFR5_O_F(VJ4TY[#b-^0Q=>cdRX2>e8GcB)EF6?/#(ULS9O6IH=[
// 8NV=<Xf]:cd84;_D_V@>HD&aE^KX=^?UTf)LfZ#C>62fddd^+9YeK9U<SO53O[E<
// 48./CE.//O_Dd)]&Wf6:\Zfe7T3Xg?8]-_<>]b=f3KL^0ReacSeP..bdaG[^8MXI
// TS0:T+QYIDc9>)^bFR02(:ag><4#aX7/AMU1gI8^5KKVS=gQVQg6Z3MeJ2P=(;\R
// 3&IIge8@T]Y5;a93a4eRYd&FTT(Q\U,_<Q&<Yc:>Y1DR-WdEN@2K9FOB[D;;K1,Q
// XHEB3Zb-KN9&\4C^LT@P&I##]<2H)L,#0,,:I&O_<FPD>=:.-O[+(dFCCEM^gXGO
// cNS+#AdB>Ra?[]PFY_<N,L0E+Y6SR^dXE,PCd#Q^3DF8?C]B9HS,1]60=?B&Z)@O
// _E6_0W=QC#J\3b3NH9Z6b>X^\,H6ZI-&6K1c,(0G2<S1F4f3^J]:,#fL+Q,:X]=9
// 3I:cH9:6b?(#()<<8ZB@Y>EXHfeTL?JRWT_fc7EacUYaE=SX6>.=#?[@X&B,R?8I
// F(I(J)Hf699@3+_XffTO:/7+<TGCN7W5H#XGD./(6@ae.:&B8]dg<-B,3#]\IBSL
// ac.eAKQ(@^+N^gF.6WADYS:],.e[JT8FfZN,57D<b2\Q_Ze5J4R<=_Ad&gY?5Rc)
// N#&^]]7[S&0Z_R&Zc-T2S1.-]a&6.V:CE@\(C/#6NMLE\<XZ;aR#0_M1/HbQ3?[G
// K4bFeCASfagD@Ye)7TTE-.2IB^^9-+g2MX51ea?06G02?Ea9@\OOAR_bBD8;]J3,
// SN?fVCQ4^G+^,.>Z<GT9UF6c[;)R<_SPGQ6D>HJ\BN<7;a8@2bS[J8eRCR?EbA;-
// S1IGVQY3/G2?cBO<./7A>Ye3X,ZT9#6N/W(GXBWbQ0[SAV:<VPOeFY&=,P+dE;<G
// ]]Y4e0>K5<W<:-EC?P&E,f8U9Lb+0/Q3WRB5Jg-6NQUY^6,4U]&bf1HAb9Y\1IO.
// ,R3SUbO50D^,^JW0.5K5.<EBQ74#V_5FOLCM^RE#/?MF.KedV<D_<RgSN)&;A9;W
// d4[V3)6C521e=[L-IC/YE/#6><<1\3</D\4/T/T)FYAO1[;geg6APeV99_DZ?DY@
// &3\WTUVDAb+e0B21eDO^^aB-KHS+C]D\KGA63W[?)MZYLd>29gUe:\N6P^HXJ,&J
// IRWPa-bCb#UU7<NPf_VX@,_<=:WFeQ>43\_E)LaYM65<1AW,&b\89WZQ-@/dXTF5
// :g(77N#O5((KYGPWf=IP>gM>Q=Ia-;):M])449e)bf.M[U+;8P8(Y+;T(^D(OaNT
// LC>NY3-A=:I#.(DQGF)184aXR@9SS>\d,,2Ha:XTVM:4TNHS9F??:KK3I@_D\IL+
// ORS4AULc,)(^(Q<VJ<fNA52-DL4/V;f56eR&BGM24=f/:4HO6NI?>KAfY6PA)Nb)
// >>()ZSc-@Xg:&47L;-.&-;?#2&_IDfU;,,X[HE5\KGRV0:egCR-U)@#1,a_((0-e
// KGeED5AV<7b)L#cIH>IFE3HEP,)ZTDTD\6OUISM^;>F0Bb:0J9W(WRQH[L#PM;Le
// ^^RN_af5;(RYcKNG[cTc[F5fEZ[IRD/#0ffH968G8gKfK#PfON0O98\;P4PA:ccZ
// SgK94A\AI(:TdS[1M;a3Jag1U)C?CXQ\C(Re8;@QW0[9;(C4c29F,d;=N,QZb11F
// -/?:&JWB/GJJ@#3S;:1<7;L9U;I06N;NQ.H7gIIL#+B&IVRd,NK.[KU7bP=/>FJ7
// [59(5BEe@Ja:PJ2(#VD\bT^YB_L&T^<@H\-bQH+/ZeA?)KFAcO^]4HKHdB)HD8:#
// ;EUa]0U9?X8OE#J_d@(N0\KVA]N<O-LP:86/W(NgG@#YB1J6D06,+b-5@8]a6fJ\
// F9f2[L3f&Z^dZe8L5f1>_FT0[S+=e4F03DUJ34-I;YR5S._>a_(?HQG5aG(,<KGN
// 6c-#D7IP#B:@D(DKA+LE#3QNOg#2)S-O__e+&9U3T_Z5d_d@N=<)BB:)K;=;9M1f
// >Q\4J>ODVAL_V5X,3D_4RQR;N(4KVM7)A9+/ZB0fKJ4,bLS1QL?g7__dVWZK+A1-
// CEO1XY-T.NM0]V,5X5@2UHL3d3TV8N(=,Cc_g]D;e=,E,=B[We?Yd[4J\EAa?Z2(
// faR?9:L#V=]._MFc@b.B3PecO8S2./>gBQQ(Y.85(bY3F>4A,W]57GKI24&Zf=:0
// g><V3D.]4Gfc9]4+QbaW7A@^FZ3<6VVPGR3NQ4C\,C^HEWR;8cd=B8/&,Q.d_-C@
// 8Cf,E&#].C7K&.fNLR.[KGg;:L.g4;ZNK-<#;:+?+K=CfBM2+:Q9g+fT]]_4D6cI
// YQPS8LG0:F:KaSa+1?8_R.IA[6CR;D,LNVX;&^&HPBdXJV[]6bbMCO\f/B=:c4,8
// #QW.PDH<)UfRge1E_C.F,Eg@Vc0-Yf21)IKWYL)Z4cE>_KNM]-L?3A7[UA8#V/5+
// N73WM_WKY^G#YWZ-A5DaI\+;6bNQ6N9R+ONF;Ca>G:7@cF/d.1M._RW6M)eVAIQB
// -IJbA^#7;Ta2A7:59Q]9WU-PTfNAR,/1c3df(,LTPARITIZc(68Fb9J?PC[PVK\(
// bC\g:=M;Q6X@9K=[/4OFN4e]_&Kg1301@K>=@:&T4R37(b^AVKA:e>_FUJ=]Yd>=
// T7M\4L7>XZ@##2,b&S.64GQ<22LSXLg,>0=)dX6C?BX.ER3>Zg5f>3HOL75A+7C[
// N,2D96C)Bb.IU6WFe_:O;Kd.VG/X7FJ^&6#K?;.>XOO=7_U<Yg7GBa1UKHfX[?a;
// 6bKP(Y7LaR7GPW3YaN^ZUed6&F(PJ++Ve++R\DBYeB+VWADRMVRH[Y8/Hc7P-NYX
// =8QHT(9Q=0QU6T)B8F8\a[,I3FS8M\PFFM_Q&4beUdSY@OgJCUJF\>+LIK0E>GdW
// 2/5FB=3Q>a:VG030:LU2A87ZV/#QCf7KE7KBa1DHLLcV@V;C+0KRg\M(Q+fBG>1,
// N3NU4NCQZ/Lf]N5)?,-ZIFBfgQ]Z])NNU5=C^-L9@#aX8A_>gL-DYH4PLY>fLP#A
// R][[6\J=+ZHUE91TWe(eKXd@JN:T,;LB[e&G8>J2ZB?#Gb]?Gg3G<[6+c)\f/dZD
// ff5\\U\b11&=A@OHbCKNIe@-5I[0_c_5=LfSTg/HUdMC9(@b[]FPe^[TX<VJ7L\H
// f=U41MWZObc-4AE11A3:O\(T6)=?3;T=X,_I&g:.(/PGKD=065d0[C>@fF)9_;Ze
// D/WMII^I^^FYN#eJ-MU\[+A0FW=Oc=.gSTdIYA.6M?\68^D58WaVM;A.B/O?SQa8
// 5RTbHTQA?T)SR#IXGG2ZKGVO9GKR@L)SB7[:RY/^&/3fVKOP.GdVK^4<C_\>EBeL
// cKJeGf#+K42YA/6b^I#=I6e[[6R@f9Y>DQcI1:-bDaQ-AD:cVbBY:.W]-A0I&ISM
// XOA7ID42daI]Q)_XQ]K11U,;.+@)<L>B@fM:;(A<f8eQdd.6&F>+MHT\T85T&g<c
// SLC+cB^EI(Ca:d_U6cfRW8CcU<[\Ae.O(gN:O35feO5=g;>b?L&BX59eOM8=&.=.
// V5N8W\=C7?aV\b<=>CE1S\5X/d4?ZgJT=1[_A]ET?a5P&.T1eQ3K<ENeB^592[E2
// RUP_2X3Nae3L4#T^H=IM^L6Lg3,.:L[]H5>\N];K.9d?(9DV=R/0<daMcB,/QNV&
// +KN2eG?8[_QWYLE-,S1@B:C^:ZSDN8cZTP0G1V)IaZ0=?/;;J+0]fF_\;.^AB6[a
// \,F]WQ2-\E&C;?SXWSTd8caW0UJ=H304X2([Fd89N8.J3QVP0>Q\)_JbFNb?=?2^
// 8D/E#cP.A/M&K&C&=9IIBN.#UaQ259\VH&3Y^,\+Q6XG/?KgV1Dd0UC/K658N[&Z
// MH;:=DY/_@HSgf&ZR>->]eCLGJ->KKC(b9N<J2;[IR<).4>#d(+S33&L?7(ZCJ;L
// -bZ;;\V#Z?F[H7SA<X22<@&(>;QM@5D_9]Z6J2KaDE.I-)TEI:(ODg5#PBceP3_A
// 9[GLAU+JLa;=XR79XeYM.da<,(IR(,A_ZRb@&<:)ZO]T6Q#bb_5;;JL2@P08X67b
// bGP]bb7_/<KT[(CH#e.NB#./PRd.HB7DX,W)?4b_1?M@a@QF2.45P+21T[9fMV-A
// 9JV01-B9f@XAK0\_92ZYdG6=8GIR/aH[TAD\<K2LCB_T:KS;V@N:TF;9/Bc1deF3
// KAZc5Va/1d_VTL.dab+@KMC+@088QfbWP,H3?4WU#a1>G1Z[]#].JH=53[d0gRXQ
// 2(\</@H0B_QGT]O1H6^]49LCbXcZ/;1_2CA\7HEV6D?O5WG=6#:D>8Ud?_(ZVg=c
// dIEH8/a8&c4IL#U4K/Y9#YU<8^G4V>WQE-]IRTBNCP\(aG-bHV&A649CLW=Y(@A?
// 8UBQAJ>4AA5Q:2PAAAUJD/1^:B:F_Q)K4S-=1=gO#;-\a_M-6dK<(,[)&,;]4C_[
// L4=&T6>GB)<#,_OL@dTb9R(G]c2=K_8QH9+A\:TFBNeHXUKV:-9Wdd40I51M/#(d
// UR&HcT^(9:.L3FPOY41)VM\LU.P>>Z-?AH920U&.N)+-5BMO6X/V9?3T/a:T4(EW
// .Q,6<OF&g4.Md<(Y.8\4g2GF2RH-:165A-LBC_a;):X^)ZSY]9Fc<?J<gNcg.37^
// Z#DFTHg[E[[J]7g/>/<>.6fU3L-SDO^P9]5\I,]M:&^J7W\ZI9?ZJG2bCPZ^]EUf
// K;NJ]+PG0b)F9F@E1Te/#R5KX,\a(D)NSDF(C&TSec@GGGT1M2:NAU^-^V=[U:#O
// IV\[=9dC1G7Ic=ENa:c+.D:&U.R?U9/D,aM<DSY9Y]VZBOFRbIKcD,94]2]LDe2[
// 5OV)>HW?FMIA@<^T^/+E8=2@<QdF4K01Hf-RJ<59&#Z1+1\JB4LV9,Vg7JT?7I5.
// 2Pd,(1;P:N<8HJ=GRE.S?Z#P=8>S[OA8R3(?C+4RcF5F<@M;6A\Z_>:\F+O:gGFW
// d/dR#g&c0EBI63@b80Y\^0X1d-Q)YQ;&R;Ad]2LM&)/T6RKc,)K5:1c[K(([+G#P
// gIeS@C)Cf<N8];,S)g5?gGTH/&J=a#LA_Hc5WR/YgeNHA#DTEP(TWW>#Ag?VJZ+T
// R#a#E2cCFgVCR8FG?_:?U+9;C95Wae4;)1RbBb;&B35[6IbG59BN;&2(WF<^>_bb
// 2/Ef?G#F[VHP:eX/f-93@g35eCOI_;Xd?//ZQP?1LNQ.1gg=UgAV(E:VL\+ZL8,F
// .BfdA8^\d@UTH/4H5#K/2dVff2KP77g)S@PY@W?M0@1a)H=IQcE>2UHCc[<fF0A;
// -VY.7=)gA,)aAVK)gEYeM^),d@ZW39NF]f5-a4g8JP<1Y5]8AG\?A-NW+SF:)(F(
// @]0Gc,UF/P5)/TaO\62W42?#/2\O@4RcIfT,bQ_NWg<AdXH,bCZc:XCX#-/fNPg;
// #_Xb4BYX)4C826HEFM1H)\P+CX=M/Z_X.TW;^5=N6c.C\YB&(.J8:PQ@2KPCYPd(
// 3@2RPV,C33Y9fX?,GVJ[MIZQ5@4BE7UQRf?E1dYT+@Y4L.=^VENK#1.eL8NXWY+d
// ZIa#Z/T8_0M+PH-,[Y_RO.8c]=83XW.6L90F#8YN8\=Af6UXM3&3bEdf\K323OAJ
// #;)8<+&cZ)=f_F]Y2V>+8M.NHbF>0^6.Kd4-BYR-.WP/[:TR;7^\Vf;V;J]UIN=J
// A43-?d/;QF8CY:=60)6,cOPFfWFZ-9-E#X)UJ9@AB-AVd:&Y7[7eCO-L3aJSHV6]
// .:BP<C(3#L]_0O?.2CAQaL@:F;SXCPGE([e_^)Aa3#0AD@UN<@1JD1]+(6NPDU8F
// ST=2,-.2.7/3.HV4g5ZQ=\XW+N7_(<[M5N?R,\-8X<3<4g(fHeBJA,F++[O?;NBR
// <0VY3Z=LHacU@e>J\;VJ?@M5&ZR2eLFJ+;H=6H7Z^#7WJSP:a_B0M^Aa/@\^?55a
// AOZ0V<_](NY2]5)E)[Fa,ARL8^<:4^L[][bD0H_#JGe:?V;>X4ROX\,\9+V_P46\
// DV01;g#O+c0I?BI7dc3KeH[9DS\]&f)VE-#.]MW>M^Dbg;8+F.=-]4Q43eZ,#S;1
// F))V>HJK;X[ZdXY[<L2X,M:gTBgM:6JDTcbb\+&@9P3PgGFVac-gbR,2V8eOO/XW
// /==Dc-1M7T;DR[A/GXOTWRe,GGGe+c[FFJA=#U30]B@UK?3C#b+c4;#:[Y4MdL9N
// L?<?^PbT;U0Q(&LcDWg7(M2\Ng([GRU/0K@IcZMV=.N?8Y_5.0E.:_<Ia:9KTR0B
// 41fBO.S6#U4D@L[5UO-:W[GP9ESaCZGZ3E)KK0N7WQ6VHfdM;3?C\#/EU/W/0CVD
// Z\^NAV.I=N.d4\V8=cO-.KD=_UQ(9[5S,g3<=VZZR5RNDcJPL6RQZRAb(@DBS;)F
// :.D,d-=D/K^29EM=):,S^BCf]_c@K;D0Xc9aN6P_)1I<+7WFQXE943deMFJIU+gP
// MO=?KVNA382FJMaUCJL_=S=XACD;G2_Uc=g^4X505?fNe:ES)P0I\-:J+a-LV>,@
// .?ff1DQTNbT++XDL;W<1_[[^ZU/_3D92>Bg:9V&&:P/W27&.#]-Icc6M,2(TKb4E
// OEGA_RF^&J&2&?4<eODe0C(CVbAac:?@U@M)Ue[Y+]GJ6O-PG;,/=##gN_Ye3H<f
// RJO>/OB6BUbK,(82TUFBUUW.g_;8UH-QE:1-5V9OMIU]Ja;c]Y56W_+_MU:TT[=:
// 6:fS1>7<<eJ\ICYUU?Q6+f&/_MZD/1+X@L)5d3Y,EYefW;KO+WRLgbECda^<N01\
// T__3TSL\W=6V@WQ#;O;bJ4?>GDd7I[BO93PHVRGD\-NT+9_\JHV32Q94O#XX7H2^
// X&QP]HW9C=V8D=D4?O0cX5L7D1?Z9b_:N4)PW?PK^SAN563VUGLK2CVLgW)NdbSD
// O?We)QL<8c?\6-<O><6NGee.<[-;eRc@]G791SVLAcR#TR6RVf7AF#\DB?c^0f>?
// ?cF;TE[C&@TM-=[bEZVV^Xbc/?Mgf:R.J^;I&J3f1_)4\YG6WVF726EeVK=ZE0,U
// 3HDB&&3(?)&91L:^fBF=cVB:@b@BY.4Zg.:W,S>(V2V-6\7C90[LY/#C&8NfC?2,
// gSP&3.NE>&7=JXISY-WZ)3ccV#3BH^,ZUg-FR=0gA];BJ-3@AK\6E,X,#3Jb;8ZE
// aP-AaNb1W@Z5QA.U2]-D-0D()b8>2+G@4@(CcX2@[R2W/PZK;4IX]SF85g\(K,TO
// JC26aZ>g-eU&\8)geaH.?AXDO]#U@[H2c:6LfCAbJF@YDI4&3P.gP9eg9=5YSXZO
// NbZG_><[McDT;bXVHZXO+F0dQH4)5^IRK366YWIGDaZdPA#J8g[H/UXV5D_9fT0O
// b,cf@XP^b6OGg.CQe._ORD]g,EE?>>_DY3EYS+G8H&6S/6_-Z1OICER<D\OFKQE:
// U+S2JFQ9NV(b\\ABUAE6[@(44H&^Kf3B8OSP=]cQR7[K-?=R#&;0FI,LEU?7&[e1
// N)&L^2OXQ,e9S#LVd_8SL8#f?=:I=WXE:)O?UEI\M@[21^N:eefI,=C[VL=#C](&
// Cg/dI781M\</O2=:A?JCMU4>E@.3f=]5#+E?e59Q-&RT4\Gec3\OOYKECSU1(Q.R
// ,#GJb9LAM[GI;,TaR97S5T;5QITNa./7CV.BQ/\^bZS.8^GSR^)E^;2L,D>b7fV9
// I#GPO,:\UB/C;EP.WbGf7@A?N+\TL&9XA]#IN+;VXC=1aY:-TN8gYU^<f>bU=aHN
// gaB3-^_c.5gLaKO]_](2SPWP5F@,6(<U5-2YgM7-S@1:&\f)EVc_+)4Ng=UJ;XQc
// EF_&D3[FJ+7BGASHUH2JG(U(5dS;VSc,)<:OGB&bfM&EP7@B,/]\[&U<;e^d_DT;
// 9S7<]N3:U2[26RIC)TKI2Yb1b3EJ]Z?&;Xd836;-KO[LcT1b95g#]Ta,3R/9?VO0
// c@\1^WgX=^Kd@cQ#e9\FSQ+Pa6ITN@4J/&\b@-S,HeT+\M(+;gUN/acE0VB_MQO?
// 5f[W_6dX\LL_4\FD2C2<f3U?<SbU_..T\MY3&CPefOf9gZA&fMEDNXE7E]_WLOZZ
// N+Nc/.#SK&f#FO1DMHV.SOTOP4>741/+g_K(#GXNOL+W&D(eLQa^JXR>)\GQ/>K2
// E<YLBA_[eV_HJN&\>ZE8E&Z+K)O5@R7VL6^4^KN<53dd:.9?Z</<8X0eXBd0;EF=
// /7>DdB#]3C3L[,N>WDR8#3KL#/bGF090+3NPf]RSXOYO&7R;\]IR0E<6gPQJZfeM
// #g8?#[)B=4IM7.=KF=V-gQK1>QRH=]g@]UO+=EH9dNS7)<D9\f<(P46A5)-\8<S]
// APUTa(g8G>;-CdQ&/-VgQQ8/b[;GOJ/GX>?GFQ]VX,93ZDT2W4W4]ZJRYVQ[YHb8
// TXNFU=3/Dg),^9WEU5C=VAN5#V^Y6VE0g1&MB)JBT2VE7+5/#W3S5GddUgWgFC68
// 2LJ1XV:OLIXTOgX?fE]4f,OG)cbHb,gF)@]9cL7HR&#^;W-9Y[gQN.93Q4==;,[4
// WSc(b::UFIM5MR(DUd])7[D(b<2&E:D5E^)e/,dMT4Tc/J45K#7K;12VHP>&>7,?
// E;).fbeZ(LR#GW]:SE3)8C<65d(P7[JWW5MJNVC6&.g:.H1Q_c0dXP11/\(a9[+=
// Se4LQd4Q/D7>.];e(LL##d4ca\,WG,2beUFbeRP,P0Q,75\)-SO9MB+)LJZ(2fO^
// 54\=@SNR2#:=<+TAX6FD]06GZd5G,,VY)D(\_.DF+aadZXY=:-Q[]\V/)LXYMBa1
// be@Ye&ffXb7]V6:LJ)S6F53Q\+I3^,[BTV\XAJf?b_N(P_cC3I6R1L0S-/6a1KH6
// .P)R<,AW1>Yb+/UW#8eG0P4/DcV]<]C4Y@GG&RbD;5f50eM-#?(<]J7--GY@@H?M
// CC26<g7^]2KV9C[RgBFDTg=4#-T5.LCKU[C&/?E;P&HC1W:c>_Fe23QI.9)/UA94
// =+[7HXSg.d,_SOVTYHb9F/NeD1/FgMF5F(6:ZZ13-O-e^@QXJ5Y)G7W>GRIR\^e>
// CR>VRcbOf2I;<cOZ6T=[A^PVPSd)2MHfB2M]d9/H?dB90&]7Cf0)7_F(gC325LP=
// >(.[?eG(eXT_8M&UYb1b3:CSH7&?]94^bAHZ?48^J[YOJQHgMBI]cKcZ>/80];U5
// -T:5+RH+a6=;B;g4MF2b6(HcS;^RR7^/V7KNR7^eH83bK2KU7(C#^LVB(@F&ag[N
// DeH(;(<.?T3-A<648;\;ODA8\QZ\ULF_-_8.TEGL?ggZ138N3>E&-6,GcT)=(;&W
// EF1ZFEZfW+7(DI=F)PEYGK2C<YQ=9^X.B3.EZF//VbX<D(3X4)(_g3&2+3L_>/=L
// H_SJ]FXaGR1@8>Y-+(;MKEXDWYI2>O#TPOM<O+S,[aWQ69L#T^IC71:LBY?bG=U[
// e9Q3+ZOO>&@=HUc4\<9&41E&Y,6\]72bF-X24;(#NR;adF<66b6@4+RN.QPcdIDR
// 8\YN460<B\9R56N7(^Q+=?1bD6#ZT\>,1ZSWWG)^+?E,gJN3d9WHN-Ndg-#5cC4#
// I@d2dE4#?I<;(X,MQQB#X-R^)3R^T9CWY=\E<,e,E+D-MDeX5Ic<A@I.::[&/6R(
// F,@K4/V_7Q-eZO?OCM.52NUD2CO8KJ930X&_I+C[S)A[>PWP-f(INg2DRBNTZY0d
// NO:>5d/HVLGd/A?==g;2^+.?b_Y3]-0KMcESR_LZ)f[<e/.5f5V1=\831;T8c^GN
// __MGCY?-);a3:PC-P2H\YePRG>bC.R-H+LX5ab#^V>\/_FQ-X6SQ@V9GTJCT;86L
// _T+2M#LT6QPbT3C^(62(X3>\-;F+N:0MeZ<-TeQKL#8BbC<\_+D+NKFE]Zd[/DdU
// +d>Kc.9VAFKH2O8D6];H>5:e7ZKUgS\L)d0KcITRDFSP3+81=PcRXU:-([1]dU1&
// />QJ]P#&V3b6;VLUYN.547ZYYfY6=<eVBGg@0[4WCd_1bDb3TGfI^7D<@ce_<<bC
// /6\#=-DJfMU\&SMQ>GPSN96+e4T?RE?\]TE:6ONA:?2]e0_gJ#YJ(YW=Z>L@0ZEL
// ^D=)/L/I(b3WLc=DT57=Ic\Ib[gF[0BG_N[+[e\<QAR#YW?N>-W,0/Dg2]TKC(IV
// Nf4?-^NZG-<)fBJE42]O._YCU4]VfF0V+;P@,=c,,GNAc@JR3?Jd/@9=S9=[,PdF
// 9X/)a7QfBA-OW&D(AgXEHD>GB]M8Wea2UVSLLBOEU709N<+P<9Qe7<;cf+dC@=-2
// JN@#SFDR]RR/V^6J5UZGO5b-;_e6IEPQR87\A_5DCF=M#B35:cd@?ecMHYC4BEG<
// &?/:&V/8b/(AHT:EQ&XZ@=X1V99MYD)8VC&:fG.9_4(=??]Ta_D9-&523H>=X,)J
// N().I?8S>^JMP#:b@=N0DWGB;g,#HOJFJ<^M_2I9/9-;E56+TAFTe#8&>LMYI8H@
// ,2=;5dXMGffFV^c&a;UB(5MO,A+J<>F(M8C)7f=9WJ;R\4YVR6b1WKEA+V=D#HCP
// 4C_G>4O3GJE42YC;9\;_0ZVMVg^=9KgcEC:3>,ES09EHIFJ2T22.5gcS=VTXA-^]
// EHN6JJXD)eO^MQ>f][_60#F:C\VKWRZ9PM,b-_+S;S3>GLdF3df]/_B?0Z:/>c&c
// #&DE<;QWECG#PNY2<>U>[(ZT:.I+?e-,&]g7)K\MPgRdZA_c:6G.gU2Q(LId+cS]
// 0X8W269LH=7;G@f=eZ5SP5L_9^dF7B;dX:aG#_9<VA0:8L@E1?5?NP8G3]H.DF5:
// GA@c\PQfUFAZQQ4aGNFG^>EfSd?a)aBB)+5,DS#gc?^a=F3XCdU)T^?[TT?@:Ic>
// ^7M.5<PUWW.Z02()WER_cKVTJ&#SV]78@09/b&=[MCKCaZK^Qcg+LL1\,Ed&6O[K
// 6g9FP]3=](f97bZ<7=cP6ONTXBSQ7\_Y=ZDg=PW5^+ANCN7QBC=14E]_Y3PL\a^+
// -#;C+WZ@57C/V6)J1^d0VdTE4-,-HGgR36e2aOb531A3H<WJ^e0:66Z)=a_)09P;
// 02SCDOL4&6L4<O7bDL_H>&NJ)PfTF);@^XKA+#<-gF+VX87F#N4Z-#9g0@46[c5R
// /HD3g\e\e>U^LUVO@Mg^>YNWf:<E40e3\e2Q4D]207;,KIXf.8,\C/1K#V7B3_<^
// fTd540dZdH<U^E>BG)E?=:W;E)\TfecY;MQ+CL-.ISO2+V9]5;G-g75AW7J46gU#
// ;I<FV=8,:TbG5[A,H:QM8XE/eg&8)BHbPP2LfD[e+/8Y2GOZeO+J+]c5\8-7QEJ:
// [8dI[_D+G\8Id=K+#:F,U#F&0GBCRCD5eZ#S&DgR?MEV->ac:)S8EWJ>XbE&C/Dg
// D,K@aM7MNG7F>/\Y)/acK01Af,+H@UL;6PA_1R-0KCSUf38T,A)15@O3>4YdCZ09
// f6N6Dbb\;&SCRRYRT>601GK1[BYE:;:H/F#C698YTW#&G_9NK]A<BZ0Qb>U9[Lb(
// X\3IR0Z9F,#_#XP_L^DK<]ANY^T,.-4U0?C(PI1VU8(&V+f#(G#@4F<6B@RQAa-g
// A^CK[N&(BAAf7HHH(&P=2/3^5ePBXS.:APDBVRR?Y.4;F\)^5_D,V^O0/a7(F?Xd
// a>#_cF:Y6)7b=B@)=C;_[-F8S]]X:>0+M6EDE8;ER8;+/ECLX754f;5Ue^N8_;&a
// 4A+2E31:(eY-S)O7Q/K6#)1<.?[M68^;>I&_RCcX:2QI/8#5/G+3-Fd-.CY.g]0P
// ++P03_C056M35.UP&9O+N6<KA<05;U#95FL-8bdOB3eY@D;=TdSO8fNW_3LJ(/S>
// 4IY(55?JQ<#=&?7CHe@e?0_.JdBN3J>eQFB9+dHWZG]a,XJFUFVNJZS2/;CK77KG
// G_2[H(ZacF]YP^@f51P9SU4<>4HF7=]EE9b1Ge0?PE1-c;<RHdP:BE0-M9PT77\4
// &3f,><B0KVb3L&TF@eQ?W\&O1]&)[-B)<(LXUR4\\I/H>6_S[D5R-?YMg280g-JI
// 6b^A1;8Z,]45J\B:E_T0cOdRA>a<?-2YG+cG\Y4TC>cDEC/0Td/<GE)^/AD<:TQ=
// LYSd<+7,1=RO30O+STgb9.A\S)>/bKJ=fRRULRX>6ZJAaP#GR_bdTb+7\P18V^<4
// [Z8g9)GaBQ]P=T(KPJ.+<Mc;(N1&&\FEHQXf_8]bSHaM7RX(ccC/BH1GHe]WN:]]
// J8+^A4bKZFU2&4+K&?;QA>:^g;Y#IY_:VGd(U0ZJ6&b#T.U(T>G0WLQ.(5;LCH/5
// 0g1;8)/Z/;5Bc[L>YUHT=&UZ/+=W)#Qb(JH=+B?2S-6fTdWe-&(?G,I[#3>02RDZ
// ]:X>GYcXQ\MU(/<\g_@(TBQgW3P,4?BN8caeOf@E-HaT\2IMRL++a^+[EFW:#>;+
// >G3)G1fFVJS<5T?S[\7@AJBU]J^IYJS_e5a;\IW9<g3E<F0CAcZ14?fJNSXDagdZ
// _CbTGQ]ZU<XL1:\N(8@J65.4W=(QZQ.-\F#8>Y7<g@#8ETS@N-0F#L2K<2,B30<I
// @=O@PIN>>IK.JZ>(D5J.Z5.[6:NH:Gc4TKD<ZS&Y^)QMS/?AFc27fcMf=Pa\]00=
// 2EbCaNa,BT1U6;?H)3+J6=+JGW0K?66]HeW1U2Y,\;bG;EU)gOWIdAL59(7F,6O#
// AcU#gCB@:OSNa]EP^V_Y?Ef649,?V@S@DdfGIX<,[bF+)bf2WN<bF93N,dCP1OUY
// g)Z<8-gT?NVPN[1QL_Fb1-;]0XLN-MSWBf<&[YcIR&T[VL\2@[)?JbLIe#O=D5W_
// J#GY,F?]<+W/&BQZX<FU0P#(aBD#3H[HB;4VT<SXLL<aQ=A1QZ)c2VQ05146VCQ5
// JQY10E&J[TYafX;:2)G_6=N>Y&dVTWGEF?53/.:2MgABB)JK9\FH(GH1:-VT/F5O
// .UA[#8-7)RAf1H)X<f.gS^7?;GNF2DHP+81/dY;(/K72Z10&K2:\:-N@7MB]Je3R
// 3+L35>fEW/1dGZW8I5)-3J0AgM>4RD(a/NEWbB8?2SNQ)8C8E;Q]_&KIG<>a==H4
// a,TO8CP-IAXAE,.X0,<TX5M(L88d>WBE]QZ@=B-\a#.a4L^Z_+3U.ARA[#b&f@@9
// E?gRYOgQ#IIa_L@&e3BNce]]c3-eeX/f..;1\C7Z]Q&b530H4VV(KYaAd-(ST;OQ
// @_?OZ1BBd\\K(We++N+@I=U^GG/L06NQ;YIa?R+,40WSU2L#XW[ILLScE@FD=6Ke
// KD=d?edS)G51gMa>9aM=4JW8J1H:9OBV9#(.Xa<@)B9I#<W.J&-6_V[IW0H=;dJg
// dHQD:fA/A=dfFXMOFF0Vc1e>H6&]DBB/I8OCZbVA/0R:NRPX=0FLZM2@e5b0/]+J
// 2T8P<G/PU3bP]RSbVRVRWF]\IA>K=<E6+fB:R)<;UeH[46,J#\E+#.)T6AJOP1Ob
// )>TA>If:,#^:ZT)(ANdTY2FPd(ELCPNV[7dX<QF6E[K+XUU_>#V6G:IQ(R)2;aGH
// ]c:J[RK&66UP/A2<#Ge[?[a?\@^Z]K6T(39ZPebK;4QC@QVgC]W^bHQ1.71KAcg[
// B[OW9WQR6QRE3XLIP_fK]F(]JJ;K>LNUCFZ;3(c#cK2[(F82/RV?(#)[HB7-^SY]
// ,?D>G)H\H(7#YDGc+A1R>G@<Hg8+G::&,WQU1MLF1aT:[Nd2_3S.3[3(XSFS]bH^
// <T_XCIeB4cXeJS6G:LE9a4#MMRGBI#aAJ.9\JFKcS/PVK;O534D-a>e3))[V,T(G
// ^U&NQ@HZIEf.bT-c0&7Wb#b7;\XgU+_cVcW]AFQB0[=;NO&.E.@(QFd(0P]L>e1U
// V3E:XR]^SO]JB[;-a1aXK+M?YX;M(4gS2AeZYWL?0f\;K\FBSa4NY\<.VPD<@RaS
// ,YZR7YU)/]L@DF)b35TDX:B^X(L)2E#4A3PGU\KdUCXBKXZ2S;+PFY/]JO>/M1[<
// R.<QRQfEJ)[RY:<>998LR;922e-OW(4(&I=HUIfgB2+IY+A^XZI4aLaK4N&+M7;]
// 8_+f]ARaeWfbPg?cbI?g-;1Z@Y+#[],XWSRS\9YDUW=+0bAB7U2A(IRMY[eF1&WZ
// a].YR<8>dYGfY/E]5gQ#I2B-?VLc#\F087(811OG@U)BRX[[DEbC?Lc;@C6;NF:9
// R#cZ<X(YDDdI332OI36]ce48V>U/_X/\L481f^+Y<g<.JTCMC+DO_F=g\4=C_-5T
// A+@O_6>Q+SGD:S_PC]5U2bb-?:2+@0ANc[V4\^;IMaD?:N;F\11XB.SU/+Y=C-7+
// gYCQH[.:FT_E9FDO9ONPU-LGUc\bU=0d73SOYC0WZfRD&FWT)aJ^OFaPX_2+=HJ1
// b+RV-A,<H#@/U5[+U]#MC1V,/Q,QM11eHNTDV5\8.8>U;<7&\1e5,1E&-8[#TA2W
// 8-M^]2.-S:=\<2@TC/RVH\-D.VY9L_PA&KF-E7DPC:aW.O9C8@<_\=#D0XUB6E?5
// +.O]b7=VGGNQ)\S94Pc/@ZReFGFaf9f&^DU^8XT]V.XCa-JA<30BbC1f2(3VQ#[C
// GQ]FU4UUF.8JSX0HE(2C<HGdea7ff^2OOdJERT.faQ9_)]ce;-R4.,=3[1=2CJI,
// gYLf]U@-(3_dIVCWC>g2BN4?][_C6[Z#aNAR-YZU20MIW\;@W1G\LR54-BJXCA@V
// =W#>6961DX[1NJ@U=Z3#.)F#VXK4(]I18(8KKgeH\)N^D\EB7fP4EEAJZ7@^HBDX
// 5c9=4TDX+XZOP7bM.^[MA?YWICP.HK?b47[(SS>J/.#[D0)7W4C8L1J(XbZdHVZ+
// #-@:G2RQE@66HFJQ2?+[GWbGPDR0<e^J[KIN8SY^cH1FfUP?N-Z];FbUbNX>@F76
// ^a6g&D4@OOUc>WP1&e.UU&X11.bUJ&Z<d)<bfe2QA_5e<2\+_MdM:1Q_e[1?6;2D
// AGDHHYZL,Q/FF_JX-KL;W3+#fJT/-_EB?:,Q[&Q?,(Q0CZ7MO;7Q-EL5HSC:W.Sf
// _VQ+3A.,IP0?e^/>,8>,X4S&:5fH6V?6P3C_LKG<2<C0.+>?Y4[&0:#4\MYW&9#b
// MGM&EeLA]C_AaPd?[Yc?ELb#MPXe9Z_/XCP+aYgP,<K6D>+GTZ#F4HYg^?,UP&W-
// Fc>VW8Z(0?M5QHIEe=#N)IW;N-CNg4_^a4=,>Y?Z0@EZZ8DXaS&8)24Jed:E\_J?
// ))F^978DR4KWY#JOB@=\5#5JB/1EZI=(P=Ia@+Y_?=(\?\-MDDcG[gV_^cB<?R-@
// 8g\\NPVOM38Y&P+BA2cc>B^J^6Nd<a8S<Ed,Ie\ZMD2/4T-bS^cGI=(E)<<]1X::
// ZBAH9FQKQK\)-5a#>cJd;Q;g+5\CNG3fWa88,gd7(VTP^4YU=E@/L-Rg_)JIEFI>
// _./--R+F_#,[H+J_C4B[6f/,=:bPTV0G&YW+bY]>gCDbAI)YUPJ]O8VHFD?NaE]Q
// =U#9)DOIX0^U(@R;<PG3R:+:gJDWNddQ8,D<6\G\2)g;ba.B]+a[7HU-F5XU0=E.
// ,XV<ZO3PEO,c[Ta_-2(^T+R;D-UW3DL1.>U1F)TT+9USN<9W<U^YVeAde#&R_KJ2
// Y_4F>18+W\:1,Ya/a9:dgNfG&/d-LCf+[=Y\XgYVf0@[03OD2^#Q9;,;X(L(c8QK
// Q[EW<a5e[O^:#G,RRP?#I;79^C:b75NJ[NKWJ4G,[VbA]W1?A^OQeUS>U(^R\6KN
// #79D9@&S/B:XFQJ;dO1P83.@0-;ZM4>/I)VcS)Q[bC(O\dNO79:KTZD_DY\?A<Oc
// QJ.V_=A5G0Q3A<J^;C5dZH&VW)@&<<5D3@f8<.b)=XP7]W3&G51e9=2K,7W1&3(e
// ZZ+H&1Lf0V.[C+22K(=Rg6GS7/(T]8(PV;.OS:8T,:bF#VJ@ME4UeXUVS=UKD+8<
// SWCOYbS:&LRBEOFeX=NL2L>PR+YD1X/BKc.OBY4B(XB,JDeF=O,TbGL2^UZ;S4;+
// )VWW.WIL;f-<,4d0Z-_F.#6a&,]VS(6BT>-D&e-S;40DUdIc)_79W5GJcU]IdVa/
// Q;]DC(4c<:H-UcT&:9[cUHQ\0eIGMASUaE)2(61bD#;9G^]b@ab.DDO&?L7;D15H
// C4&e[c0,<94(+>@W:)WNcN1;]XEK(X-@F)FAC^UV>>VNU#=Qe5DFd0f_g4b&F;a>
// 47ZSgOZK#=M_a^?9X1UK6JBfa^bQ@08/5,JE8(C/<L;+E46aFW;FX<b<XfSN5==2
// X(Bf?<=Qf005Ea3MF1,9=7P=9D2Y#/,>e2IHWeS7GD8V?M;Tb#HaO-P7O0+DR(VJ
// W3C11OB8@PUa/?35L9VfT>TA=S?<TOLV:2(@PKc:1A@\9Ng;_/LXf?N2<H#<aV_#
// Z_B[67)=Mb^GL1(ecMH1[CgW@W\0OgHea>;AR_Aa;QI8Fa&eZ+[NE@PWg-;fR81a
// Rb8ET#PL<QB(be9+YF<MZY(>fdH<.NE13D<_<eY,(3<PNSe(A^W]g[L9.1SE1F_b
// Ga]KKcb;3^&)#T9^/?gLUY=aXWZSF:WFVOeO07F50I:6gf)8eIMLFcY5Hd@=M6,C
// ,#fe3[[<DY\9@IePG9T2L(-=[>PCH&V6[6Da2UP-ZEY_ZK,:eN1@K#[&d6d,R9(d
// e7OHRf?AW>ISH^LWM(,L9BAC\TId56@BK3AdH&&-TT^/W]>^LM+-HT:5;=WE:&d7
// b-4/-./T;-ZI>W(2=I]eQd0g,Q=&0I?W=LOW<#Vg>XFBWV_CIJLg3]3IGXEe1C53
// EdC+K(=^&??PQWV1CE.d^B;+;=:-WCeE]c/XgV1,EdX7Za<Q8AgKFX3GL3ABW0[)
// cQ[YJ-J<Z4UU>W0gW\Vd;V?1)M@98#,OQ@J#:E:6TONQXTH+D=@[1:LEY[GJ0@+K
// -0aH0[/-Z9Q@L=YH+V<.9@2C&SW&(U,b.R-_=+=c>6Ob(8d6+gW/Hf6&/[21_]7Z
// 6f,#5UO/B)ZL/=ZHIC?GeMB0ZG(0H&dfefZVUF.747FX[ZTNBD/#K/G#[8B=+7U+
// K)Z-5Vb7QBT?DH#Q7K_<80-@;X:g^_+J]-3HLfd3G0[c.W&_-fQ55g,dS+_dL]+W
// >0[/YOA;NNT1D0b0YTHZ:>Xe,9LC7OOE(FES8d8;Xc1._aU3OeQa;R8W<IBC[acc
// g5GeF/5HCNR,GCCF]7J>8)1)Y>Fe?TBA2S19BL?6&P3J-5^_fd7d#b3&M?=_7+UM
// )BLKO,W^&Q^=17RQ1;fTe1-3g9#JM^TU1#GcVFa(A2U/TV</H^cD<Z=&7R-PCG3c
// C<1LA15.L/D4/&)6^A)=aeBCVV]Ud3;9e_OA,M\,1dEbLC?d_Jd>A.4,450_:9d[
// .:TdJU\bL&e+07>E^QgTOLS;Y#EU+@NNg)NI8bOQ/#+2UJYJ#8WT.X(S;UN_)5QJ
// #N1/SV;&0DcceFUTLfR1F056>;SO/&EF.1BDZW.TDWT>=UNJBI/?ZB=2[[Y12J[S
// 0:UN]Zf/Z&)Z^8F(NT;9eY^KM^;F,(cNbWA2Mb5TI+S2+\4\+=/<24C;fW(RK^A^
// 3+.;-5PJG24,AM6fZ_&5T)5W)g&Q0LN+P)>FMX6+V\-?@)eVUV(@L[J.JS^Q1XS@
// (W4YG58R8VUd[3c7F&FMB=Y/^/)_/F]^OU\C;/7AaMA;V].dEP6M.]f)b?K;bD1[
// D&LR-a2I0WGa&S?#(&)737^:GP6QJVTL#B8:.\gGDLH(1HI<#bA(&T0IO&DCcLTf
// JfO>BJ73IbP?I-N+P[bNU90(#^O/W#]^OWHF;G6X.TgC\:96:1PJ1bA#T]YH^)5Y
// D[)\fOg.A:@E3=3T\C3F1=A_fb/F+[99,Y1&6G]M/\1<NC;GFb+NZJ+5fD)YEE^a
// /4/?G7P.&6#IPU1-5UYJ,1K1(?EacY:M?,K/@[>83#cY8RB?GB6=M8W/Ge/QW.@5
// O:/cMM#[G_J1T&9cUG&L5C8G?ZIcVI-_4P/HH@cd:JF<g11\d+>6DA=6N2P_/WAC
// +RUdEL-T<1Y^[2:3RCe=[S:bf,A(=T.E82HU?.d5U<;c\[dHB1JYd:c:LXPcUROP
// AcIT[4)gM@)RDHCbe9agfB,)Hfa?X7JMM8G\b@(Q>f/R=T]A7LB#@\3D7UE7eH6F
// ()KA/KX/6GW(+^8GRbMP[G+dC:_XZ.CUaPf\O<1KL-I>WRfLI0SC#_<>ZK0)GS(A
// GXB]NSfb^db]f#_bX0_K4=2](N.WNX)MB,FE,gL7X7/BbDUF)ePB&)A0d0#eCAM&
// eRGZ9>T+IRS;CGAdLJNAcb[gU8AE2gB^Hc]&&Y:9BUK#;L0,#RR]K4?bHO>?YT^@
// \g:3>OB_Q;5E-^P4Ta#DF.0M8B:>\2.P^T\\e:7?d0.&TN<aCK;ET?ZcY@6QG+=T
// :4_F7<]6S<;&66,=[>.D,U-9-XB.&f&2>U_HL,K\F9B01#\TNNB\#KA&2+I36CWC
// <4?GW1+8O+N6>V0W1[-)A>f.WI=R\)=C-K]OBEeC;N^A3dIS6;7V,eVL3N4B:8Z7
// :\]/=f,(H94DFEe8QBBG?(K<.F1:ZZB=BKNZR)HS+3:.U.Q>R3?5VN(L?+(5,Hg5
// DJEN46g=C+1V(a??H\cE#U]?)6COD>4Y,U6FS5APIO:9]M=];QFI3KaE5)1-dKTY
// &7C@\^fL3bMDPIYL;NFQ2#0UKXTMT-(?KRd8A/&V1GcY=VW[aBX^(QBdS>/K24&)
// O39V2[RMILb]-a=]@#&X<=0I7J;N6,BYWQ(aU:8[F;&N582#T(9#P)I7PgaG:Z_F
// 9YFfc>]9Z/MZ-]f.[;5R\XR<g)=7;V&@KcFc4?GfTVF<NOKL8+TJVCL#[JB+8T.5
// #]8<R@[XE:^&T-+)cWJ2BR0[^C=f><AX&4fS4#[5\a]ZJ+E=,:89).L)W6c9bN?]
// .(K]9X5,2NYK#F5Tag3?5+>3XMJ4R<Y3<CM\YG8bRCI][8))?c]OU\5H>EM&Mb<e
// F8g9PN:I-<M&1=#Z>KCAP>Ra5bdM[4^eWJ488W0=>_Tfbf3HW,44[Y7_;<54#:M:
// RSAReY9:[DRH=<WP4/YQLV8[82J9AeL[]B)[b=52TDSH_)&:Z4LE@gAdT;=).DGD
// 3d;7.X\/=Y0\N;ZOb:>NBZ;<.:G8;CTQKK(8WU4gA8feV+P;6SGOQ2M?3+G&aAUc
// .MHeD.>+^<30^TPWQVaVRP;f[9)+)Z,F;O=1T^I/f,?aceAJGQaHXUHRVHFY<]6b
// _3:8M0;RXQB3=F,XKCUU[8+4J7XM@TKB\CH)T/I9SL,.4f.e4gf-Ae:JOCVP1WKF
// M\@=G;caWY2H6A.5OVG7S:.IAfUD?c)>)>KLHd2d_ZdSBXFS+,eSeD[=e>H@Ug&Y
// VI)P?]&B/]D;\G;J;9)c2ZO6bMJbK1fgJVP3]RI9_M=(RCBc:;N++#8A\P3PT6W4
// I[#H6[J7GBeV(A3T:e=?d6,N^,(@FD:Db>/^9-b5(BDgV,5:\T5Kb<5Lg:T_MaPT
// >KB&4/U&cDE8E<D?L&D?@+S[]1N@DZ]@S=DOaORd5N9Y6c<:Fe9f.QH9(3<.SLF7
// B+HAK>eR,.U\)PINRP)H4Y(>=)0;T(HH(OY=Aa]3,QDgC)<+RCb+TU(F@9EY\A?K
// @^,f<R<;Me9YVH&WW&=BF/\CCK3EYY#)^L9EC?RK:>B@PaJc?@_&_UWK9T[UAA<N
// dE^=IQKAaYge.TM)]2acYCY6[YWT5<6W4\#d\QD>\B>UU1cXcM@L:I_>.@bUO4C;
// ]K,aaONZAG>@;PT[41UO@J@)2fMW@-.CUM@R\Ma))Bb1Y?=dJ;]PFHg/8BVP:]<5
// f3Fb7aW5PAZB0PVPN(U&9&LP:CUNeVQa7;+=C,[3W#V8@BJ^(_&/8\.+QX&ZEVIf
// I)-&@AXN82>7Y>/HGZbUA]-B?JDEDaYFNC2GVA9W_fU6D]Z>Rb@E<AC<H_PUWG03
// .WPX2Q.4YSS(\S=d;<g6KL0Z>^OgR36)52<JAIH4J]\dXKG8Bf[dC>8/=9)Ac]H8
// Wb=Q&LB)&38gSJFSdR9d\OWe\A.PWQR5E]?&SSYRS6W(47^0DT++8SR^g-7/N:KR
// 2I<=_dbNU9Jc8e)+,]^\4Q6U1QYf^aX@-IB=[IB62\U,W#gb895UVd:8bb;H6:@G
// BWKS3RVE?L\Cb2F>1..aeP>,dZg-(SWH]CQ)bXgGd5HZ7cO[,/_@AZVU],\C]O+J
// YO4>Z_F^I2/cfK1[:2-=)A01)0@>D[VO/f\gK82PP)X+#>,I58ZgI=0VNJGYM+Xg
// We])T(HgV9]EV)L=b:MZ0OE+?Cf7-F)1L6,PTHJSNL>]g2/?c<]U)6<#?a(/<M?[
// WfTLGX^a[cHf.aB6e]gH][ebD_DNA,?=S(ObD74@\e:GA,APC+G&)d+:G#e>Z0C2
// g#.9K9._\J9=&^WIAZYYS9ME;E9.6A9ORF7.TRU]T_c-=,7V]SM/#N:KI_AXMU(/
// e_?Wg&/g:Z(FQP6S67[YD[Z6?&MdH<Ic:=G(26)>U/XU9;+4?f\BME((COKg1YL&
// .dP^4=,3.ISZJdPPK/\B:V2#5FM==eB?ORP7X0.#\^)c/H+7TF9VLKTLCWVW)/EN
// <6=7[[3dedZ<(FaYX.T)X]C62TJJ:E7B^A@]a^\9-<4>95.S:P<Dcb,&M.9&Z[I8
// 4C[1:6T526Rg&X2Q0QGaZUG]GL=5V/P3SSH9U0\U;H-Me9?/_;,Xe.gD:gFgLZ_:
// FSPR;g-QH_9PS7H:@_N,Y7=d50R]_#dZE5HFA,Fd@KVVU(?(30=0gAe@SB-#)]^>
// /?U&TZ,.I+31,^_d#(bcdO>@K?D27+GH(f/G4d<R=W@JG.U0TI/W7Q]Ce_GH]?Tg
// 4Y-R+[[XQ\5<.X<7./?#87C=CeMb7C9a5^YTgU3\cfX^/5e?I/G_E7S&+HIbF&0\
// TU8[/7NV^NO1_U7&I:DF,4Z(LKf4=RN1^L11<NGA@OVGUX):NIQ3>XWD]#G&eP3Z
// Z.;?YO>=a:83Y^M@eL#HV1Vd:LN#9)64WIBQfCe?RKZgG4HBTW6UD(LF7L\-b-YN
// [FNfOOJA7,&>JKHE&1K?9<ca5L2cNJFN\TgTX(V(-d\L/FL-9JYZ;4EO7..G7,_f
// 9=IIVQO&PHE1\=A&7,=\-bSPJ?a]?A4&[,S[#HWB2@N8#[7A[[PPOcXDY/1a4KNX
// 2JCbTYM&/Nd;aF--V4B&dYN/RH4-,ZTBU@?e-+=K+&(?[B>-D+E&HId)&/Z0(](#
// NG3AAXI[>+1#JML)Vf#&cf<90dS0f^;f6)9XDYg79W-G<e.=76A3&eV45O=K+7;]
// 3M=+:D>Y2T7?#NDAQaM-^2>T;A[1&5?)gJ@N8)&CdS^cWOd\BR6C.WHI]\#\d+.R
// =RXRgZg_bUO:,6CL?VJ\UYFT59A5IRcRR&TFJ6_1Eb2XG[C,]c.SN0(&d4OSA.94
// @HgfVQ&YV#@_VJARW<1AJV283^gX:=W\U@N08@Y()F5aSI(C\B41KBQ4J&PAZ6P3
// d/I9=N>/MST>\.V5,E/G58eIR?I_GXBY]fd\O8S325J&3B60U?K6HJc,0&bE:ST[
// 4dS;IESD(9DZ=KG+C8;LQQ4d7O(Sf=UEG:FKG;A>XZ\_&AYcTXDO.Q[Dd9N0WfH5
// e=/67YOI=X2U.bA-N49eWX/ICa6E1&&B2,I@)Ub;LG1BF7P5Wa\MKbbM&)7E]SK#
// .DFUX@(Af<YDHX0M8;98@.QC&_KQ;Yb?BY[D01I1=6c->aF,O588f<0@4PF4<PK4
// ^/#@R3edC2EdU\0H5H;;]gBUX0UAZe?[<?1ReBWR4cT\YQGbM-),DdEe<)EQS=>R
// LS>Jd8ZA8@:g<@1JF4_Q@CE8#J#MA?B^VDLE[>JX)LNBAB?#V-PA>_OPC5:YQIRO
// @MP4-Y3<0))]/-Sb3=#WeD9G0V::=5aGeBKW6OcYXOf:T.]^_&9gV^1\MLI4TK<D
// FbAa\Ma7V??^CDA@R1GMUL])7DRNA729D@\eG11?AQDBHSFOKOcKTSbOc6_>0U43
// 7FUY/Z?,X.0](d]:1S\=Q[N5@Xc>\:6C^f,AC[[WX+J56cJ,3\g;NDYW^7#-VJ7a
// WWVUWSSUA8)cTD^TQY__0aW7,C,/KRcbA2L:YPXHbffJ9eZcW<W:R-]-IeCFR,.<
// UXT>AS-8.]\:Ng3\f[+=B19EgQC/.-;Sg?8+N7<85/D=L@)Z(Kg5SbNd>+EUF_Eg
// WEf<f7HH>N&4)O.74<5E:>DI0,L+@#@Jb&_0==KcBORM7BXbcMIM<@_fKB>=e(F8
// b_DR7HU1/@-RPf0?6Qa[K@S>83\2UO]QRcg(DbQGSIdd#GKGA2))@G);@[[_JK<7
// 53T/H-<P-]Z6H8,VY/XbAd.Z2BfA-A+dME4R[454##HW00>gT-YbB(O^#UOZ?#\D
// TZ]U&8T^09\R-Y0D1V:=9LNdH\1?DWT-2+KL3QZY?]FEQ^XWQR.KgU\<JLN9T(HA
// 7SO?T#=D<3/&2R:ZU:C[:6XPQ-^a?6VG+(gaT(&JO_CA)O:FL]\1])-:Yc?f?J=]
// [4VF0R)IL:C3XRPB)De_:M8=ER0I:U3T&,9<#(D@0?.]3_9;d.#APb_S_C3BTeAe
// O:UcZL3dA-bTUgUP0:RR>,Fc2e#c6=A7XbI>Tbd7JRG:;aCRK_NWA,SJ<P-Q-dX?
// S4-RE#63UISHYN-\4YHa9(OJEA1E<I-S1^D:V:c^HGL_<fFL>TcfgLX:XE]9RR?<
// 7FNaE587c-P@U^8SC^5R)G/a=dCOVGD>FHIS&3[SM3EHfL#Q,8FV27GUeBKD(442
// 6aBO_(9([Q7>_OaK.e2M8E.10J#^,#1D[WIg-AIY^)MS&3gCfT^&XRP&0Rc&_1A4
// &#b2CXKga-;b^O=M<57=V.aG_^PCET(FJJFF6MSG2.;?2dX0eIgd;RY,ANSeNc,K
// 1TR?9N5T=c(NK+QSWAN4CdY,e.UFO\SEPJ@#>ZQ9Pd>AbBJ_1=TULgN;:8fR02IR
// <1c\[&IUX(+>1Z1=>M^8NR^&RRWe^]0AHa-FB2bWI#)X4^HJg1,DJUQ\82])P.CF
// 3)[R&2>2O(3R8\)Fbd>dNbWP4]/WJ::)7?<J0&-+d5WP<,6.f(N-:N&I,9fR/#d2
// T(A)<R.B@(M[[@NN]F,6AJF_O^S9;07[W9K(T4QQLS;[Z20Y?=aaLRP66N;G2R61
// Z(IVdaC\Q\S4&@?-72TSQ]8LI:D#;@DZ1M25dQB)^QMcJZCM9UOe1;9YWWI^XI>f
// 54OT,D14V=30E]dYEZIDAKg/F:0Y[UUWULS(^AX.cUe_.PW/AWabZXX7&cP<P4^2
// Q4>OLJdOBCIfT;94eaaf1N8,D/A8bQMb1-+XZ.eYVR&(YB-2.7&D+8<D6V66KbH7
// ]f)]6HeOP0Df\&ON9M4E#)Z.V-M3S.V,BD_;]@>-d(1^aP[=Y25]GQSB&RZ2^<EV
// JP@IK\).1/;^NDJeVDbggA2b_+TD8[X8e?7[_F1A;M]E=B-:<WBFe+XfaVaPM1FS
// WK[\#PeAM\4#Z7?E>@THgFeNb>OT79]>6:Zb[2,R]?7U(Ra2)+.CE-L83(&cP.C;
// aWGLPJRMbRN;U)FI^N]e3O2L2SfNaJ0(^PSSQUHMS;EbQ1WKH?f34WbKIY/)K9OZ
// I57>Z^^@5RHU^R74,_Z)-AX1aR2[NJ?g63(5NBENOZ_^[IF6HX^D-1gV4XSA?:ea
// dGF,O&[J=Z[:;@S(SZVSNWe6DLN1-b0@N-R.YQNPJ0OC_cN8AU#]N<07__,)gDV3
// JNf<([ZcO^Y0UYO3&1@),QU)e_X>\Q5=Zf4gYgG@gJ&2&.3Z<+?^4e_J6[MWH4?#
// B3P8VRY;)&Q=R_#3RHgKJ,JI0Q15<K>KcdMM#=14W@W(ZO)A(LFBV^_9GGMG3HAF
// ];&O@YWJ7?D:ZZIEAFS[ZAW:@.Id3#PNZWcQX@S;3;B6R-UQ11VZBcg]5^[O>6Q,
// DM5&/U(KIYCX:6d]Q)MIP;\7a0Z@/Tg5ZOS1g06(7&#79[T.[&5HV[d0/([<:O\d
// +[-RB.V//7M[7Z4RX>\DU.9:<W1Ic11;;6__AV[N1V,OO(f9QbYN3?beIP+I\&,U
// 0HO>^4N.gAWd6VZ0G?7[W_a9b9g[@M#e.AF,(.YZWN?VJ,aRNSXMH&<Gg1BN\3^)
// QF/0-eS[RdE9de4EbA-P.<(+Q.+fBX<UJZ&B/0@3>aBYAES=XDO\ITGQBG<6Y3,6
// PP3+VT_8^/Q@X)@7,2_2)67aabS)[5+-ScKEK/7XS58B^65/=HN&G)0]_XH:SD,N
// IR#R#SC&<#Mb#]e,1SDKKD0Bb00C6XUW@ZS<fcP)Oa_&d(D02^A,ZaZFL<\D3#])
// eGg:8:Mc>,Jg\&W)7g@@&If^)Wgb-]#(2Hg1R^Rc<&EgW1(8VTGMMRN1aF.-&-Fd
// +2IF_USQ8.0aTO>gc0F:53>18DA)ODbZaXcbF+RA,a+@@dXBA,A?TKJS6I9H5,/W
// 89JJPF?S;I@I_\MgPe_@5UEN]P;0g9651I2L/TKGgPGR^C1eCW\<=R-.D>ZO@c#g
// bJb>3A[IV+(V+f1RbE]\aMbD^3Ee#+1BYf^97Qd>KU3ADJN7W>M7PPQB[]UD8/;G
// Y+6=6<>;8f+]c#3LILGgd[=J]1D;?<86PQSYL2Lf9CP5YCFdX,J8B8f,/4/]\U1d
// EgP_U2G_gNdU[+bY)ZfYa3QYgL&JYTaHZP/CS2J>/K-.<A]YF/)aMD(L5\/,+4PN
// ?T4[+,bfC=g73X?Ac5]g;0gYE3].M;\C&(F/R0588\b)a>_)-QV1FS>gYd\CE:82
// E):[fE2ZQHN2HY>YOO+f1YZ;5PX?7)Q?ML9D>T[4.b73ZUO0.cP1?N3V7_c6fJV.
// XaWB;N\gWDa>#X#;OWYB@9RMN;T\O?:bG(,\@&KbR-b>F<^H)bUa0QM:=I>BQJ#W
// C;QW6ZH7(GQY1fN.?-3\>DJ/-ST:\\=GL^\YUe]GAW@9H_YBD7NBc-?HT659YT;:
// 9?KMS?Q52gTdA.5[F<S#W\bMK(AXfeD=U@[J?T@@>FVgf\^IW76YJS^K(&<\@06J
// _K-\2A:O/RRY:aQ?SU;DR4]Ic73[NWV,e0?C?HH@YK1Ofa1Q<6^UJC#He,.<^)UO
// \SU)/=)g#:dD-6@-YH/b34,e?+[9Xe?O25F],bQFRJfZW2CO-6V:2D(TQC.UVX#^
// ed9#Mf_EV(134aG:Y,K.;U;&5dC,&R,1(L:B+/>J)eS2[V(cU/,ANQe=^JM[KNB&
// \4HB52L2^6e76+gRJ/VMR-D4J>,RUJW9FPND\DBESa--DC)O/_+,QD\SF\-.Q[WJ
// -WFY;^CbFUG#PY]3U<^0<R<+G=EC+HR0bf\43]@)@6#5GT:2KUP:BB=ETG63b^PK
// QF&FJbOS=8^..T7._H[[E=@?</.6>F2c/^G_;>6)QPLHMO9)^TDcF9]bg.[K&BQ(
// LDBK2)e5@9#c7.be[Y.32.3A(Oc\H_MCXdaZT,fLRY2]M#8g/[/VbXL:OSIA1_88
// E_,(HYXS&D((UV3AF&EV(,C\+]+=)b4ZfSLe=)B[P#AHf^/1&/4(J)b8.-]6P625
// \dWPc@RO[WA=0cWLd).4cc;?FL:^CO04RGICE4)@1XTI&H.;C6L]-GUD/#e1N,7?
// acVdSUGFC#GY9<E9EKNOE9GYVHdQCQFHN623-:Z..?RCf<J_5B4KK>5=N3J8U9L+
// 6]@,X:-^E?Q#FfcGcWf=9eJ_]Q&)_1H(SbT\]g1cKFO#<19P_;VfVZd\=eAc?-@E
// )_8bU+A,#I-37?._Z\XRY0(NaI;dgZY?Z90aUcH(8Y^S)D9F&,.9RM#g7BEB07QM
// =).S>4\WgFR@?9W4+_KEP_6SU.1YgQD#QIG2Q@Ie+GMZHGR.ggG&<JWe11CV(X5;
// 6..DH:Ea@KSVMQV;(_#H+e79(F2AN2Y6BH2SH84?ae36SXX<+Vc_W(.H1Y>R=(74
// MRd27_7_RE3<C32/R1)=:aC.9YP]_NJ<^X.^S,Ka@e9b)>K9Q]8#bCI52H=AM@JQ
// 14;(7,7&D6/ad5V6\SccSZF+&_+WBI^OGe21<[JY&.f[&/R#YEI;[X72P]EB7A1E
// R;+2+5Wg^.IbeU4g9?.3MdT7AT0S#-?YL6dZ8g1AG[9PP]HS?K/LE\/KMHC,Jc99
// -?MY;J-5\Z+8JZ-E9cb7K4Sc2\SX^^&FX\#LI+[[>97\WKbeQZg6X8MOX,F)Pg,0
// ]Je2T3cLL&Q0EMG^SAgC+4;(,bVZ_/=fNT/0?R2DQ/2+?^G(J2a:5I(L?PBN\9ED
// 4Q#MKb)O9_X@/LPYGZTV)7PBNU^^7S_1\9[;CVb?DR@+?df.MG,9dd95g4OFJ+Ff
// ,H:-+7+(WDFXb@&SB?g<7]LSbWUg/_Ce9_UVT1FRJ?#A,XaV,RH.,120K[<^RHY[
// =BdH\Vc&J>QBC8O(:cBJC[TG1=;,<3\[2P#,X=0VR6&d_].;FII9C,?eg2/M1V08
// =cKOY7BFHP(<f9&;;,,F;e:TJ3([&]DU3+_4,[cDBgL_0(ec9W,Cg[6/I0_3ZR<R
// N9d9][1&A79a9AL.NFBR(K&2d=J1P]];0?I_22-UY>VeY5(VI#Y_;eXA.YGD0+[Z
// .))7]OgdXLWK2&AJ,32;TaW^KK0&Ka_H6]=N&d@#&#BSI;HFSdR\<].RLELIOVTV
// geB4f:fc9dTN,<\(>#AJQILKJ[C8feKY=^@+;IY?EQ7_(fMgBfBQ36PM,43(B]^F
// VBA]R+D(=&D,M2>IHF-2:P^Pg(VbAg&Jc8F2,Kg/^WTC=.36RIJ/?fS3@TSL[PVc
// L3:I[e1W]HL#PC(PCA/c6];8_BdEgJ(RFTZ&<9(&[-dg/IS+4c_>#/f0[66Y_[a<
// _LQbeR+bLL2Q7XOe6#6-H-G8fC65;/L41V&>ffROSdG(=b8L&9<WA8QO4>(RBc\A
// ,3V+4YCH68;Q.3P-&0ODZd4.>Q/(O=BN[Z:NV)U;4P#;dD9C1b@O5f+N5M<P5M4R
// 5#3g^0I311558@7&\]1[Uc^d/BH1>ObOL/0gVeE7e[gZ8=.9\#7@D4F#BN-XS3\F
// Q,)\2&:aB96@F&:;];a5F82BDOE(3@8BJ]e)B@6#5-f&Qd>I[NPMBFUU-FQK)eL?
// 7gC;P).(1d,_0:@W@fE65S33f^I@Vb5J/X_L,YV<EHAYX-6e=bAd:e&D_=3/U.QO
// ZdL=U;=B1bb/GeYe0aV#OMS?O7cfH?eF>OF_ZRN<4f^-H+VLTX8BEI4KK^]A\I;,
// TP?g<M8FB7^,(2AG?aV[ZZ7=TGG+V+CZ-#&O.d]aYa/8)V>N-1ZAVG<OZC5XIQ-e
// UI)A&OVY)8UN/C@YJZ3Tf8dL-C,_=U+T+\0^N>^c2/bNHMVcG_CZU_bd4T]^RYP-
// [a9=1.86LXe7a]><@ZEI<>f<e5&;AU4@JQY.46e9SL<+G^(I@RWc@-LHCbXWEeM#
// Mg0.(4CIF4JX+:aTaJX0KQEP7[N@[5ZOAO9X;d)N#?5A21f_B[EZ_=35XD]JDI7@
// :La(XN9EP)+)E7WU9d(C4O;]=b)8YaH6fG+5OU>5P7E7Y)=AG<)XXA2^&\A^M&>O
// ?ZN+X(.O>\N:D=\/a9eb[PV?:^RL/W4Ke<.2O\WS-X+V@++;WRUa7Ede:4Z;E^4_
// ;<0[::,/_ge1eb(5/-?GM]dKH_IXRMJ(=f1AH6][Y5L&5M[#84[g]T&]/<R0<X;f
// \cgAS_=C01HUH1R&eO447EZ8Hc,;&d)OHG+g]8_7/Q#IR9[Og\Z:gZC4=>XJgH.=
// SP-<A8?TCX4(FeC;=\aUgF:B+cQ=M/J^eSOaY:g24@f9&Q5:C_I0#./g=VV^.2fM
// 4KLMdcS:4+EUdcb^6508cJb\(-4@)[cA]Y0>2::Qe@VD,0(AA57#7A,3ba[Q+;MX
// _?I\=;F#0@,_?&TWD?3J5ZOFb4VI\8JUb[0?^PGEO<=:L0A^(@RO?[6PDV]EgAG>
// dU>]U82(;WRJbSO^[NPc<;\;+=XXg62gfZ,MMVI5dQcRA6B=]LSJ?:H\M^JM_F+W
// (H)K]F=dV/Q7;YT-AOMc=59Y19EC,;)86@8SbOYHNDe-AHDQ/^5,.UeY2;.e;8Z4
// R?Q<MX4,<EgdGKKCUQU&IMYaG+/]WBEMLc]W+A7[ec=VFcUb/K6eH-<-)V9ND)YR
// Y8#.NOYKC44YH>JS4B9D_4Y387gf5B-H>EI]^+A;&9T\4[eXGJ@[(B)0H2L9RbT<
// YMZ8^4:X5PLgEZRL??(/?4FD0M)0\fFZ=:YP09@47ZZ_9MXFT[>C8U(?>OVS3G(F
// I++#C,\fL:9.g<G]V/O.6#\?+Y86Z9bO?MS&-5/EDC4O:g?(R2+B,;.T0WI<)GCS
// F=Y[Q?ZK[G&AL?b\_^f<Af&T7C;>34O[bdAHG#aGPcg)1gbg1BH7Mg9@bKU(PMab
// 1J,G(W#L]V[,BdVRWLVRdG]&7VbMR2((e6.e]D7_?7TWaf][L9S<BJ#cMR6B^DG&
// 9WX[4ZGC>c8aLfBVdc5NC-=J#3S0_b0^:BEX]J5_+&O8GU4;]B8Kc<N<fKOQAF^f
// F5696F8.N_9;>Gb00AM7_XJ@&76S#HHCX<?e;dbbS56g<P@WUK263NHO#QP3W(TD
// ?<E05.2EGb/;KN/_Z,T)-b/]YOdTZB0e]&aGS17)6.Sf\PTW>eWZA2/-,1ab@N2D
// >=OFDFfQ63FbLILYa[H,/[O9S^8Jc],^Y8D;+GB?54_]c59HA0+M/O6N#O8KW-g/
// XL4dRd/@A>6\5T-AHLFDaYN9(e)D->;[E#T[8e]Y2eUZR1VAVXMJZL:a(0A8C0^I
// .&53EM_,4C#V5YKMH1SGHQ?:Y2/ZYHT<1T3A7FS7?a.//#:7HM1IX(bF]75^HW#:
// 6TE(^CY^^V-<F2#+8?&>E-YS,0&AX87SOA\GQ@=0(X=+b-8bOA1NY>5PMSE5f<&?
// 5,TI)#[4MgJd>]EX:>@+@4,Bb3OfE6;?bb9c/U?>+TaTJf^)2cPJ-dO-YY22dZ3d
// ]X;O/67He4Y4^R-8?J:2M:D8ER1f=Y:UK+XIVS.GC1Ce57f1])@fJS>(Ma1L\ME0
// W;&&2^f[NGBHgP]HD8A3EGED++@EgMEX-:G04)<O?UNES3_9<D];#:HaDc([&VU=
// ?M-?Y0Ob.A78E1>HVWCT18Z?Q^-1@L\dO-#dMG_=[PO,FW_Fag@_I.dG5a5U72C1
// /d6)A=3^ZfZ4IA2YH/XC/2W[d+)TVKCFH-/JVNZ\M6(5275OQ_#B[M>\g)54PMO9
// 4bcg[_e+eRg>YLL?cY>fG7&?eLIMb;OB^:2ad-2WT@ZZWdd&BHF)1e6P>QfOT?/[
// RO3^=c05FIG/+_?256g-MM_T6ZeSNC2>^Y&XT\d:]c<S0J43MS2?S[\;TCE&V[_Q
// ?F&DTCT0?6Q[9.PJI/T:4b\&6GH8]ScCP\R8[(fHOcd+:XW_S>eN1?RNgFEg&O>@
// CXYB]I#_:N[S;4g^AU&Pf+eO,a(8/U&BG:(J:1&FKV1@gFaWI2RO\Ng_YQ#GN<@+
// J\7:V_9/WL,8NCDVAN9UJ&8-^)CVM8=#+JJ1/7N;C]96JR<Bd;(^8K28Na0A^R+I
// /Y4/dG==JeW;-[3ZK-e<E(Q8NcY12RC@<,UgE\L\&TA5a>L):N]/EM//;B]GWLg/
// 0Q:=Y;)>cVZ>(RG#^+f\e-MVM^<YF>]T5S=4Oc(_FE?>ZX.PPV?Ob.)O9@+UX.b+
// KD9X9>PHBQ.38@C=2G6@MV\WT^HV>1[3>gd\X32&-d<\&^a.b\UFe+2:=DZ:<((X
// /;#SXM>G]_#W<#/fEHe/2SG24;L\MKF3&QJa\TCTGQZ_WBaQf9QAd\0;cMf.<]96
// VLH<-F7^LEAfH_83WLQ2NYg=5+QD#CG3Z#&F.3@_(^U?&DJ^+(GW)V6)dIW,Nb:3
// .;?(9,(2-/\35PFQ8]OeTd]IC?+5UM0=g6G,]0RScS;g\1A[@Uc33YFTH-RHV&H:
// _G-L_94[:+_+&^P^J-D0OYX6aN7a]-)OUe.O?;[WZ?C@P_J=TJQN)IS3S&-1>=K&
// =;;#9>@S]KGH]ZaeNQOXM3dSZ@g;[ScY7BP1Wa)+1-+S)<eV4E=2E7&T_E8.YVBP
// (;eP[R-NTUPE=4YL<.bC7\A=,2=H<:dI;e6Y]-)bLQ]=Z;2P;WJZ=A1AB#GVUZ9Y
// <HH#..?3)Q<RfR<E/@Eg>[FbF0DQA1dQSa(8;\McZ;RE9HYU)&?>7>V.[8;4IfO5
// M^Q.Q<8cb@_)EdW=#FIg@51.SUUQKIKB3@4E3QG(\>8[<Vg0JXQNB.782:&-U-\I
// PK@\B@VJf5)]2TT-.332OQ=-\WH?P_R\U]NV-?=B?8#[28XH<:?SBMD;Q9Ce6g.;
// \)Y==1:J198UL4ZME.96dNZX8JSG(7fQd3.9.7^RMGST=9J:8YF>YREM^@O#,N,W
// [8Iba::UI^-2-gTbD@U#PB8_\bE(IZL8T/;ee);8:(.J,e+2MI84@4K<6=M)P+I3
// #K]D8VAb4CM&@dU.:]O&a_1g[If3^OKc[&.RB:\Hg5@\OWV^G.eE(#JZM(9>_b>?
// cN23NUZN)TH#9(Y:gYgbH[)NRVN/Dcb9S=V[DT1Y0-H8-TL4,:^c@0I2MfcI^e&0
// Y^@=MFUSEHP<HWYc10B,_<G^cb5S@4Y7O)g76W5BW7):?ITa5#[A#SfO-C&dQKX6
// ABIQ(BWD[LE,5-@K;DX0ff8OFQ+LL<\^M)30U[b.^8f?3:?_B9XQ:R<-\]AQ2&ab
// +;JgPM[^(<M\_::<F[.5TW39\Oc_=c6##QAHV(Y;gQZR8^4\7M866aDAKAF4U7L:
// F(:2bbJ5E:QZLA>R)ffA_77a1J7.F3BO,UeIWDK+U8/699^8X4A1?)E=8E75ddGV
// Z&c(X=,Y]V>dNK?Q5_fg<@d(XYa2g371-B+GaA\TUNV;3RETdL9CIRg4ORaS_;;L
// b,+dJ/P8+<c>-7N,gVQ=J6S2U>_FJ=T][gV1@/G#WMJLZ_Y@3,#/Vg)f=2XHWaVR
// df,<AF^?7[=H=WUR_(+=b3UO[?VQN(#1@d0UDIWIf9CcI31FR>KbQWaK7@QEC,U]
// 5:7KgPPKEFR:XA05F-J3DL/&gff>AYVSDTSU8)FV59;gJB8#:\1SC_XADS90M<6P
// D@/A[c&T;W?Y2;[.9KTN&7K@+SX/5gfUWXX(bC+_SgG5.]<<0QQa<O&N@<<MZIJN
// ,4GL).UVZ(NYXKE_YPgY[4CW+b?>6+\ZLGG5gM+:6]Q26OQ0a.QEe&aUO0B+N5be
// &3c^^NJ6^(bDG_7K[=X^7)0FQ2DMBgZb31?Qb(==-E(.MOPG06ZUa8Vdd/.=PK1H
// YQC3@5L)U5P\&d]3#6AG6G\<);+LPHcTUIC\Gc<Ne@9f;QeTe5:b:&bOTW5.-eWK
// I&TQe<GGXfZLW97\VZA.X)5-eIe(NF+ZJ,_8C4[J7FDCRV5NS@VM^A>8,FHII3)\
// 11-,RV#]JITZ=^@4T#JWYOAQAMFG#,0DZ2eO:[b,KWI0_Mc:K2\Qb+fC<+;YGd<f
// 0,\-/cHPF^R;]Z5eR/#8fLV583@<R>ULVJ7\L.0a\bZ^OS)HdOBg50BSV\2(cVK+
// gW(@WWRF#]&7g3BS_[M4:f5^<7HU[cBS_dgC[F0?OIJ.-8;e8/EBX[/FBU;,:Pg7
// Hc5,CGU.9GGdJCW?1RfgVMNIN),?dId3Bb#3?XA+Rc#Ld>D,[6\GFK.?B9U@CB[H
// DVIY3=eY5F2S)Q3DP&4aALQS#Z._)Oa0P?&^Y&VI/7@,3N.R]^_H(2;Y+7:#)3)D
// KJ;bOES5U@]+a#e\JM]<2BQIP^LX,a5aZBff#2OKQ79+d@-V6K&M^X0&_^D<Ug6X
// 1&A3\T8f?.)B;.gCTd,ddO,V:ea3+G=U,N2V3#QcVe.J;J5[J6;?VN_,ae+Z58Wg
// gCYLM[USF0WWg47\HQa:#1W>_R>2Fe;a[0,S7L[_?Q41>a>aX+WN?,MH^e,V]Q1X
// @EbLS^1eK6Ae990Kf>,Jg8Pb2G;1:+aCOFLC97gZOZ@1XCbOD-G_?b@+;52HHP??
// WUCP&43EYSX_(UK:P\(dg74Q5[?0Ze;0EQC:cIVM2F3NHTGMCDb5TG:AZGN,K?Kc
// cKQ^5K:g>ccfSX_;3Tg#/4(E/QWc,4O>9PVf6e/Z50;,Z8:bbD),=&Uc?&6(48W9
// (8?IS8IM_KA,Y.2-TANeR_/>0(-Y_]+_+[+L/fH4.e#7[MOG)dPYO^X3Y#5)NLX(
// (R)/__>bER58,D__F+=/@+#.D4OEG+e=5f8e\<DP;cO0]_P[MYI<YRd::_3YSSf/
// =#/((<#SM//NS<b7^3LH;<?BH\T9#>4cJ?G5]O)81V01&dUgKAGQ]P20#Kgb[KfF
// )Y<eOeaO2KF7[SJM3d57Ue6I?a0D30YNf;)7MMWd^Ca]aNI@+;J?TbTI:>[)ecWf
// \##,VdAK[UDX6^K/aW0.<D+U)IT_?df5cE@3cVW44#7+)X6IP?K,1[\+9CZCR_7;
// \JVPFA=0V8WRF4D7<Og0.5\L/:L/N5J\+Ag(F))ISX[T5I2/([L_FX@B0b+,3BE8
// KEU]3f3#&S1Yg+]FJ3AO+9>Oc9Z3Veaee+LR9c_9=.QPECWgM0HdN\YZ<TFUD0B_
// dZ7&J:e:OKY@LdZNW\F_?7;.A2^bC(8<SWQ650R>Z-gWUMP.RJeTPV6GJU8?=,&,
// 80+3;[+#C2NS5f(S_;#&?4WbTB7M_gSgB5=KSPYaH@ITIGL)G8J8]^49IWWYU+^A
// bGP3d#_G&\ZT784aOK_P?W1Y/GX@=9+OLe;W=0FZ,Y(0A8cR,cWHPOEaFVE#TBBQ
// SK?_J?S2K1[bA#1X.3OK?+ec-9R7.W&P\c&7TTUdM-dBP+a=+-\P5-DX5K.6&UFg
// b6>&1EY#X@B&bSg((>,gd62TU:YG?0JAOLeYDW;0+H8eKaDQ_:V,J,(dE\[M^]Mc
// c/\d]RFaNf\Z)B6DAbBLXd//#&Q9RcBE9IE8\O-R-QR_KQbT(1S>;aD_=c,NM;O8
// _O]2U3C&fe1K[I@:gI6U),B8QHJ0O)/-_G55N_HW64<KNBZ>4U.8P:?,#,LLcXK\
// IP\Q)S_bJ56\70COa9&U9CZ=6.4K;MIG,EW,E#7D9JKb5]60M]0f(H^:8ZU24]_[
// WILOYMb5.eDGVOPUCSb2,U(&;SWU0E(O8NAZ-2FSVFX;\TI3N\+ABc(,.GYET_6J
// PY;d>C\-[4,dK/?D:[:K:\bDFOHY<dDWLeeCE]O7/eeZD)X-cS)M8Nb;DN_4BF^@
// I=g9P:889B\,,9[7Q2^SJT(S[?871Z\UVI^\Y8,_E_;.)#@8UeX.<J8(I+e77T6:
// M31a1NXS&>R959.K]^]GK1F7)e7bd^BO_.4]]d)K,4MD(c@4L,731I60C2WXe6aR
// SUUR=G_#JA;W>@1HMaJc,E0QG44,[I32K[M+37&7PcOD.a,]#[U5Z:HY48b@dY)Z
// c]=?QP53Q,N(U;c-MNS+#Z@;NO>9Cgc\91ef/[Q<RV]#B&]_/C6^da3+L+?0QW8_
// ),LZI5:J7ISC^[/Kc<1<8NPN-S^I29H25<V4bDVeg2Z[BW(M6Z46IXQ/,5:;+baC
// DT[R,G;)[527&ZAa+V^B)cADVe=]:_9<2L<Oe)Z#69RK;0XH&3GbU=G]AXY(MDGW
// 6[/Gf3L7@D=b+Gg[FXRBL)#4,V\YBU:3LR@29OY9?fT/B21Qb\EUBYK[;PF0I8+5
// LM^A0[9>M6Tf894ID;MY@.IJFf7O.LE.g/ZdR;.P8DU^U^/FbfJO<39e0MXL>.Lg
// MT7Y2]K_;g9fZA_/:AW[/VI@,\/[<_LbH1;NMS]5SE00--?.DY/AOT1f0:MS[B4Z
// 0,6GfC(cN,dMX0(&=b2NOC@)9;TS>:C(EILNT_L.+1)LC=W#DRHR=,C#1P+=4V^[
// E4gE?d&,9C7?EbC-&F4ecY]dZ.6D?g3LLT\5-=85ed@)B4;6.SUYA(2:eYS]U+CO
// @>-)TWI#6[21HL7N\#0I./(R7KG8=RS]^P=-W1B7IE(a,;>K-1<9(Uc;A1XBe\++
// d3M]WT9[+BVQ=8,J(J\E=:7<NB.P>P5@)^2BK)Q-]46=QX#J.LOe2:E-:4G6TC84
// DdR[S2)O,J[[O9&]5)ZT9ECI77)4KJRF9\_Me:R8&,YKFS44I1&LT\)bK,6=.?^Z
// Q_/A[8H7-YZS;??LV.?UXNZ9?UNV34YMbRb_e+X/d+OGb72P80<]:(-3E_dffL9W
// ]->dgPCPg@Gb^ASf?M.9Fg3X9:8E3fCJ\E9A8KG:M5KTH2IEIL1DagA?N&&X9[<X
// feLLK,2O]d5TP5[^E:UDC73eRED(7c-Cb(QY=Z9</eO(MI2P8Lf@N?7ZLA=c,4--
// A3d:ZZSR>6Pf0^DWKf>Y>FK3&?T)2ga08GZARO++/C?VV4O2?.PgNSH0;a/(>FP/
// (KL;U)B4Y;4]Y&TB8>^W(Y8>@L8C93gL)5RC]]G7&6U]FG=HQGFLP/:-T6]/\&CM
// ?MHZ##\c:?X^cP6dW+VL.R&d5^TOE(OHEV1Xb#W)b3BbF)FP_);MFVJ_X=OC2_T#
// f_49O7&D-6\MbM+C\]>:-UVGg]881XA=I39(TM5B07LDQ@Q@f6@)#<W-fLJa8)&O
// 1U2(IdXC/g:JP)XW+?@QLb,OADW5W3O=MED_=T:)0030VK-X:f^c(_FM7d3N#gOc
// 1-NBc8I>b_PT9FBARTO-8gSf[^8P3P:&<QGGNP5/IJ[+UI,6J#RWU8g>Q\/0:\[F
// ZIXKOV\(7VDVe^E#I^]?eU56[_TENX<OVFV+0,M7T.M[(/I@?eV0=KgX#gL\f,@I
// +J+DO78L<SJ?[Rc8Q<NR.-3RHW&fRZR(.77<IWgUG=E(gZ4GS.Y_[,dC8GXSK)Sb
// [)BDNbNU2(X-3UE=K?\VF/;=C\&IfS(YETeT+9[<e:=ZJ_#_g@2dAZIB0JDfXcdS
// BdHS3VF142_dHc\8-d.B65+gW6/#g_6;cRK3;[EeS?&Lbd,[<EQaYY<;:[d8&/A#
// PgK[KKDFfUI<,PZ>A2:[2#7C0]SSc)O6?Te@d\(QDQIJe9X6,,Y(GK?N]4@FF_(L
// +BT@G.9PMAb2HS^0W,QR3,#8V6/Z@W6f(8NH4U0D,5WQ_.P\3Vg1U22d#&\E+JGa
// GV>LGEC8SFXA[6B/5VaU1&7.Z35]??7.J&#C.IYGe\23UO6d/#[,)7KMdb>)ZbZE
// J..f\K2I-@VG3;a:Raf;#4;G4RT^:a7W6Ga/C-6QVE(g]:L;IN]dHUV.D=4K(6(1
// #\3IX6T(2e/19Zga6]<J#MeH;dREUf3/B)@JS20O]4<+Y#6M&V@<GBWdQJ)Z9_73
// A9IEHU_c6#(@aG=DCNPaeF-OHQOdU9Z&394CR0:U(<.I3?b3?G,(,&WBO\KDO=f/
// c?(BV]dK\8IB/\-8A&a_WSV7S:eS2^O=5R2&O,eC;/:9XMWPVV.-BHK<aVddOQ1-
// #TB^U\FK,cIF9UT;@2Fdf#_3.^WY^)eeUS01U()d<6RIX;<C8HOT;2Fg65+e?#^F
// ,\E6aQ)8ME+ZF3H-HB#Yd@INQU;T:.SVLH<Eg,0CF_#c/8L0?.aT94L0V&T>:b1(
// f5EPIEUOP&S)6S0SaKF3&6[Za<6[D(.PX>U,/4&1,/490>MMcfCC_9[g9)DFgQ:C
// X[F:X;K;_Y@]KKFYeOfW:?^;@9.GQR6IN7@I)_dI:\fWK0V-aJXg\1>B3]^&#I<5
// U/5>Wf<RG4\C@Q>,18W;g)AaRRB\JYaQ5/H/K6=THbf(EJ:UV0b(23bD17Y&8c^^
// W@b5C]6RAHSKN)U&@[ZE@CeQV:fFX7OY^bRP8g)geMTRa_&)ec2S)@6aID].9JOe
// d@AN<8(QOY=K.a6JY9BCY:1E8W@AA[X(:<d?_@8POL5FWUfg3NcH#4\fRH:=;=d]
// >;Hg6)J.Ua95;&C&I0L&&cZ&.;]AOY@E]-M^N;.6<R&\_2-^.(-74JNOS.RLJ9[1
// Y2e>)X\Y(.EMd@TdBS)H_+.B]SH(6?>P.(AY_Df5\>0)ETQg?d-C7X9J3c(]E&3)
// b7CE5^=WgH>4]1VQdb0Q=SI@63cI2[\93ED/C[2E\#SG_V[^FJ=)5]&2:X[,<4<\
// \WA-d[6DX.V2+gX#00RMS^8OERC\E8J0HT_@P9?ZN7F8()+M3<9D.@G^eRe27^YL
// c9S?1NZ>eW(MQ-V-Z\(><.L=1Z#e]^g,dP-)\Vdfa&712<7I=O]V0Z:Ec7M_G&9Y
// XSAgJ[,Wd(Ld0QVA&IDIHGG(g[eQ1eXROa/CC\Y:.;cYf#1[(BaQ5g;R+JHeb9@b
// U,.PW>LE@C:9&Ve?VUPf[DdOOSV]aaf7LIJZ#W2aM0JC1D4.aNO,MCBDbaK>8B;9
// /7?06Wa:R48N2#T+CJ.20QS8=F+W)?U5JKPL?;c5#X:B:J^dg7?EFA<T5d1U.V>d
// 7[4IN/MCX]aF6XH1KM>Z?b4d_-N4.Og6W@\OQ@Z[-3.g_BgDKdL=OA^AMDYV5LZG
// \eS]UUKSEB[L=][^GF4@S>/WKCJF+0da(27N=^)aP29>ag:O98Q4H^UK02I5VZ73
// Hab+c_<@_7NLX_@IaJITMa;cU-5=#J)3,B#A,G>[3>25J;NZ(4>a62aLO,@Q\8Oc
// B=W?^&;[P]:Q.aUN(,/dI.IRW;7,VA??=_(VKV=]Pe[-Pc=77X,I7>QXaCf>R^C6
// ?F:;E=&;(R).MAQ21D,RLJ)f&ZM>DH\YE\7X0O&HRYbb\@4+Z2,BO,e&+=gCMH[6
// ##1\8.CS)@1g1g=gJMD>6=V3[eB]7bUD2.-c2I6RB=;RRN422>80[<HB=V1(OeSP
// \Q^71d-XeZWXe4,fdf;c(SEZCaE9f2>+,dJ=I6_ZZf&b5L74ZC0a;dbW350#&:EL
// ^SZA7+;g4UD3;H7N/FefW),bb?gQYDc4,1gAI=54,OcS)L^L/C.9c0]U<I(5MQ#B
// QgbC<FE@2IFO<TE-:V;EfJ2CLNEW:K?BNM98<KK(10aP2aQf[Z)>P@-P;JNHB+_T
// 7PONHA&@DBeF9G-,0<7I_3@TU7(+RJTCR9AV0B6)3IeeE<=XAKJHcM;EK5N<Z@YM
// @7@1?]5J@4Pc4e^CJ?=>56:HHag5=b+I6\;M:ZcI;gVe]XF?WZYa:Tf@&dF3UR0a
// =W#^U(XBDV-QHfJ^\_eG]M(/:XSY;.X;.I@P0^)-K\F+Q.fT[,>SE5D(,SC;L_gK
// Ta>TFX>L.<HV_Y.A7)&)WL_Y<OJH[O6_R>P-B/)O<@-&:(Ee:BM8I\<AJW_<?\0W
// A=F-<0&PfLI=d>]CJK4E4RG?S<TgFX:R(VQT:?J1R:(]K&&:^12[T,\CH]JEX)6B
// L,<RD(,D-K7QC5Y)402#G.feD5,J2U=Y#LT8+R].A/0G=)<O.4DLZ)e=1YYW7/F[
// XYX[D8>(8[/b@<N#H0J,eeYMI2/+CYCOUNE-\&MR\YC09FV7+F2=+J/+JGJVVSSJ
// #[?CJY?T_)8>IVR,a7)8GV5G@(PQ=;B93[F]6;/1WX)]0+TNYPg-Q9A@d9&NAgH&
// gWbL1POIU,U(H.FKWL:##.Ve\3cY(2Z4D+1@cHUI15RV/O,CQ7/)B66[/e;NRaQT
// PZZW/Pe:aIc6AOP?+),QIIYI(7S:HIL2Z+Z^cg=>dI((U73CEJX,T8_@-bGBb#,C
// PB=LC=QI?1/Y:=BfPA4#IDU2EV[=_)IIA/.gY>QeFD,B@W)48,2S]1^^QcWKG)(U
// <<RLF8@SaD]cecO:8e(HaK1<KFL9069/3N^[/8bE?,)D4&_F2G35NL>BVLII4Aa0
// QN1KW?#@EQAaRaDe?W?.@BHJO^KGPXG+VYe9?[HL((_-a,37-f:b9Hd@TLRM=@+d
// 0Df\@?>+4ULEd#bP9ZgegF+S2_S?FJUUIaN+[fdS=12[3)D8,^+eXG<)4EMA?e]E
// MVR7F/(6g6Y/dHWdQeS,BD=GF):A&#B?W<Og/WDY9f.A;:9E3>^=Og5/_9;E9LHV
// (&[2dU:_KHA;JR9.C#YMU5JaBGad6L,cE(JB;)AV2FdS#ZHgX)QI[/8BME&8P5=I
// 4NcPF1R[2;;\3geIPG+RF(/8V_M;098eAS6-dO#KW)D8(&W[]P;Dc[bDN45/:KF:
// SU?+2HFO#;e=f2_9D4cA99dLN6[#7F#[X\CaH9>RHX[K,5M8&L0/BG)0]YG(WUN3
// 0/)D[J@.fb?.I/3P^WcgJ6U)7>--UP-8JPKF>R?_E5BD3)9OP#/]Jg5f)^bQ^DU>
// NGG1>Sa#]C(LD<@FOR:WHL)PK)2MAR5OX/dPfLYO519];#N#71W?#NL:7C,R=b-3
// 9,+Ad9IJ)=30E52ZUEBOc-/1FPFgWF?]&R<G5[L[bc]UcXLZZffTa6QO3<ZL3<.W
// IXMV)VP:>ZL&4<_QHKS9Q0D/>IK?d(#-Y9UO1I)BB93RBU=HV<f[=1JII<N/Y9bD
// cBDEW>7/EgOXNMa/LQIN<EV&97JQLdWQ;a&X]eB1G#SQ:X(b==/M.Va&ae7Q^Bcc
// ,f2^ET.4[[I2R39U,]fO,S[UIZK#[\RQIcE>O9LM,7?LBK4&;^R&7Yf;JSJ.D>5_
// dT:MBTKcDG(@C)9ZEXO2^R,E2G3+N/OE]TO&ebK,[^U:C<SSZD?\g\@fgc7#)L21
// _4TQe-8V;>DL8=:&U68OQ]36F++<[:d.0;V60NNPFKe(Ug67e3&5Xb>J4KA[fL3<
// DO<)ARH5#9TPN7Z_Xc^B.=3Z.Sca=be7?>-.9C#52-]54L+^6]P7DC1+Yf/7M.C8
// 4OX5;V@.6-REQO]8e56RI[HbUXRe0CVCb]dbRW+R\++<]Pg>@3,LR7&?80[5L\/&
// R^JK0cT&Hf]JE80+BOXEBTW)A0T@/?Q92K2:CID?d2IOUW-fN0f\YRV#[c7(PP8f
// f0#;H#2:=PV]/Q=P&=YT,[H#AEE);0aO_]J?=a^1.OCH)Y\/GPQV/=782]EDM\gc
// TYe#NLC2^d)&5=^G:Q<b/B900JdDRf(,;W:,5ZGE8E/J8CG)_D[M8]5@</#ae#]:
// D.)48&)Y]6:.9G(b]SX0;H/.;31#^@[QIO&;G34.]Y<WKF)IgM2cR?O11LY=+(Aa
// b>aZad584A@bS;\11OSUf7S=4X<^^M4S+>P7EbP4LME].fGTKM#5.Y0+2YD\QD(1
// )e0)RP??T77&DFe>^_GcC+1)M?SXT+RbNWF\#[22DHR+?G.3X-]<0<Z:5FcZcb_6
// ^)\@e2:&ZWCWWCAS_eWR-IU1=b87V9aK.GC_;CU=8OBDSY=8fC(5:Q1eUN^;(K2B
// Cb879BL&O4-gI-Z;R8KSSZO.1_Q/JUO.<\fY+7c3;]AB.(=SP8P#NYD9<)0aGg&d
// @-=UNIF7Y,Z@/b;N\O_BEHC)P./Ygg]b7G0D514[XW._::b@4gdG_W=G]Y<M<TEV
// 1bL?CeeQ7c79=.CQ-I4?_J&LDZe]6-3Y166f6M)0W;IK>E2Y>5=Ya^CXC;N3&Y;/
// ALHF&HF/9Q,B[dRR(F4_aAVHB<.HI5TR=)5>SJbgZa6-eF+_?WU#,R0f6;C2EO&A
// R)H#[R-<S.CKTO>-9VQJ&Beg69]3CELbKUe8C7>6[d_Z<VJPWC6e\5,WK;<-27&S
// MC<YM,GD1VaEV64NGb6]-B53NC3M:O5]ff1,]5)I#R+9dVc_)CFI#6?>V<GTcW<V
// C:ZV&+6;:C9^5V=HBL_]aZM@?;Cb6cIKT;H5#,^8:T[Vb63gU^d)SaF9eKXLA:0V
// K>2LcL=36:H\HaREK+#KE:(_ELaIT[9(FM)F[IK&TQM,ZWFZ4MC86T8LIWWKM1<S
// NFgAb2)-(c#B6KaE1d:W\ObR/_AV@M>A?;UZB<(a=6+FTW)4VMe+3Q9TE/9^7Y<;
// I0+N-I2-);c:9D^9I]?12eSM:fQN2;D0f+gO+0f)-X/9L[8P4WW3J,Y]agb>31f[
// ZHc..=Ga=@(3;DS<gQDN3#LZTPf+a]BgFX<g1ZcU/X;[.AJGA<Z\3_:b8bO:VV]@
// 8DMU.c@W=.&#>\.JgFE2+&/U^H9;TYWIDW;9]9I?AY<>L9A_\Y&=PZfW5_HC_^5V
// Q5-6PZc+SMI&ZTF>L(YV7<VXF?0AK8Fc&e6f<K>3YA[_2RBQ]G/#d[P8?IP-/c6P
// >(.]J.&@(6)W#HOb.9DGKa;g@BeOLSc(&f<@0N\9VFOa(ZaI]HK(_K4H,+?8(:5<
// 4);\?CQ(2BI)IP]_\@A6bF)6SO3PeVbMa^dOZ)#D82M;0feU),J6b-D7Ie:8&?(M
// fUE\5QS=Ug8\)WM4S4)=Q0gMZSbH@.)I\7aPb;FSU?3dbf--T:SF?K.[0_dBUcCV
// URVI6ZDXVBERWI[\IB2._))cfSb:[5UO_;<^NJH/D7Q]:a9B3M,-/)Te-Rd;3PgZ
// NDAYX5ee4gFFK25]=&bI+?9+PgBaS+H,,S5,\5fb?7Z0eLbYdfMVKL.WW(IXD\ZU
// ^,Gca_OPH>S0XLKI8J=-+AC^2V)^bO],I^bB1GH/H^:=ZHI-UU]5+#X&5-\0eV5B
// BG,X\(KN1_/2NADH-U3HLbZdI(M&<1@_f1g1JV.M7(0RE]N:5GQ#Zd(?eU^Rc\>S
// /::f94LWU)<LS/(Mc7<,@Y+XO&4I[+H#=H6<[19^NbbUK+6JDC+KYE3B7=fD0N\K
// X9C^_.YB#]F/C[B89(TRXMK_4Z6+)D4UBQ<d97GAT3@(HA?3=((Z?\0Bc7>@-DK2
// A8-OM>,c&.>ARZ0<MIFN9I-I[Y+S?HaODM/Rg<#TV3SRC)AQT^=cW3N&?XEgU#@D
// .X5\C7782cCMX5\#1B[0P79bVT.6V<a69fCH]\f9OT<E=adH,E4+31d]:/<P.4]f
// 53aV3L^06=c8BaJS?;[,@\Kc/^+BPWg2cS.9WJGV]Y,NLP1b8f5_Ae.TR8C#@X(I
// 6\>[+6139;ecS)/-(CB7H6&;?GFS(DbUc+L\ab/Bc@]Ce9S(<PR?GQcCcL,J8c=.
// +/,_e)-Ra@E-I?O>d=3L)GDS7.M0J_10a>77E2B]C#8e:7CBV/FU;B8b,E>,#5PB
// L4CL?:/UN&?LZd2cRD&HBAaeY@YY9O2B8=#N\@/3(b7H)aF.4K]2==LF3?]<5:L6
// BKQ&2_^f6LNPSB#UD.0PdR00&a:MO25/H7B27a1O=eO^4XUNO;\2aCQ7QK#NFY,N
// YfQ#@A\>W:FcER3F^BfV;5M^&WQ0TPb?E,&_N&VafNBEacX1PU+/^f>OBeYD>B\D
// MYP23(JgCF)EL3gS+L5_g\+\A(fPRXR&<\Ag7Jf>;HDSSTN\>VF?ZI<(#M5_K^R.
// 2=8Z1DC2:DL/.SZ_Q]VBR=U06eD6_<[LC6f1A-;R+#Nb1G0\5.aTaV+(?F@/D-fe
// N9ZK8)g?gVDe]1<e?Qa)=#W]M==/(MZ6^NPU@adZK9#KJ5gGKX\@K]eO8<JfTbR:
// M]bJ]f\/72EL0T3,M6[6Z[YaBAC<;+--ga8(DQ^d3c\,Q8-UE3AY:BHfK?V]0E,&
// (Z-5NQcOBOFF[FRbd+28UG07J#Z#cfV\T>Y;.1O0JH?Mg&0X=FMG0=T;&@,b[aV2
// XCW1FaJ:)GZ8ZeCBI61KDCJHH+2FE^.GPZ=,2>MGEa--WdR5SbE4,(6E&4#.=QM/
// H7QG^/?WL9f^-L9aCT7[#\cIAK.O[OFKRH&P7R>7b5;aBe;EYg]LH\W[RKPRXSI+
// ?VYe&@X&RU2C>Sb8@;g;JG?dYf]N3=PT_W9f&D^)7UBT=NN&BB?_3[?GJ<,)#]<7
// DK#6<aU/5R)D^78VXNca@A9dd/,NbG=aTac@LC03H1a]gLg)RNVK:KdcA.-d^gWU
// Dd1J&Qb\[--[&XE?HdB5I3P282,GG788C5904eY025VM>XBZOfMH/b:,UZcaQDe(
// 3Mb@H.Ig=D2-[d;:eR9a.2d&/AAZ1N9U+>M=2I][0-8RX+XMV8A[G^)@3g@@NDCE
// d1B_B<_5PcD6e9.UW0g2<B?aQd4\DFZ5FeN_],CQKB-gcT7L[cDKZ=?B]2PQ&HTK
// P7f@?GM0RXB>8P,_?I+5LJ.WS9P@).P.DU@OH@BSc<fS[(g[KSa(803f:#I?2dF\
// 9,LAP(:.@WD,VK=-&gL.cS/P;0THe-_9Mb2f:#DFM[5O).&>cdVX284V>db95ceV
// T::S.dV+(RaN,KQCf8CMM5O\JcWU3;P527\<L8C[3X2G,.3>U=K<AI0ESBg[ZH8>
// 2U#1e5.E]0DR)FGVD55]?)[/_8EJf+c-L=OYMPK#VA@>JS^B;a<8U9X=_#gJ8?;F
// N;84,&AU\<_QIC;eWQc=B8.EC#;F.41c(e(+\AD8Y/2ad1^A#Kd#?+OR\_3H)2Q\
// TV5E7.0EB;L5caS_8Oa/02[H>P/Y4WR&2gbR2OVH(T=4V]?<_b48/9\.WS.V)g9O
// )^Z,F[S#C<A/CabaA,d7#AC7K;.Wc8M^XCO<C9U(/c8W29e\MWa7P.#O]7VCR]W0
// =M4_3(?K,UUZFBX@WC>@NN->YE(CYRU2PdeId+TCQT)Z5Bf8&VDd08HE]b5POYc]
// /EQV3?Y;@gbc.3.dIR7b>O91c6b]PL[Z7Tg4L-eV\J15bccSTBYb8e6)RB.N6YO0
// -0f&;H)3@V^QXAc=SA^E7_0XD+gON,#E+A>6T1HbA-)IAT4X^0F[/9f&<VH5&T3/
// PVMZ03(b-g>/1a&^PV^EA54\:@0P-d^A>N--C?-H3)@A5G6(]5SF-EP(Xe:+1TIR
// ETW3BO:;BV+4HJ#K<WQee.9HWR:?=MgLacN7F];#^RBW<@,UgSWEb[9)efLM+aW9
// <E4M_TTYLC[cPSc;2S4[Q4^E<[;650a2JH^7H.cR@4U9)UE93]D,[D+,81f>agL)
// B>UC^=Y9+)a0Yce.gDG?cA7R#:Dd)]1L:QT7>=<@TC]]ZLMHJGKbg>44CT>fI8Jb
// ()DdU4PFC]AS>-:H=+HCW]2GED;)FBdKEDD7+.X3a,8)bD&-QH_6@O6S#HU?WZYV
// FCcAf9UPb]&_c8O;3I]g2Eg]JOH@SN>aJ:SA98.:P.:d.4#VKSXI&,KFR:0WWP)Q
// SXQ?:W_7+4)_1]0(3+95RO[S,1Y(-=3\a-.W3I1CQgYdX77f5^5=XX(&W-<@9^b[
// FF6:=Q99bg.g6VP^JJ&)BUc]P_BIYM^e^:V_PY]]&83]?/96&PSg\(Y\g?EWd3/1
// FfV4P0/]Cca-<8EE;^]TKEG]6fN?X:8LX\Zc<1_1R=-_7HU2?N<41+[0<72@FdV)
// &SL>Y>dbV_g7F^Aa)T,b(O#b6SX[(A^Q-NI<@#)5_GPAMROJ3LL,b:(2?3bQ]S8T
// ,12L96&UPKLL0C>9CHC[NFTGU5F30/5X03PU466MS4aOX7.R8(faf_8<53=O[5\<
// =3=4=MOK/.Q+?D<T/75V6#I&D@UZJF,b#;SN9C]\QZO2BKc\N)H5dPU3e4cTS\+R
// OfGPB_#\QIMd_(c2>fIg3=a&<4^HJ#+;Jg<C.M@;RK+L;2E.B-FF96f@7X7>[0/^
// 1ef/_fHOOW=5<I2R?7+)/-1/,:dHPS#_GEKDX[QMOUQ6KE?F,/G@:VQZAT[LK2@;
// /ePc2Q]B.H=N+SM\8?A:Aa=<@>E:7+O<T.g;F-5]O=^6A-Pa9ZS3O:TJZJ)2L,:F
// ^2=A_A4C@+\Z#8b:^I?MHbKWYF8QUY5ce]0[P-=YB[8\Xf7^>R9AB:H])30EfP)>
// GEC>.1KP/NaIHC1G(8^?XdZ#P:O(a5C3MS9ERZ&1EYOM>B8W/EPZCdGf6bP]]_d1
// @^:Z/YA.A:#.5ZLO2T&WE0JEA86FO4a(LBCe_U7@E=\8?:I\?>X4T-ND;D47PQRb
// VK>f(OP+7=DRV@6<eFABZUW\?;U?c],3-SN;C14O>,[ZaR[^MS+Ec6WOK?Z[SeGb
// DSBd/g9@7cT9I^,_gYcM+G-EWCZ@P-LSEW^I6^P@gYBYKW,P:a.,OKP98XE?@4P=
// ?Yg#O2DdXbBcPKPY8A]fdYM3C/]TP?=5R52.Z/R-d6H=cKPJ3O;PM<5_B.(IKD2:
// G=aIPB;,C90^Df6,PbW5,?dW7g3<:I+&V#_-K6QV8C?&a\(I=f4SR]6X++@=@DGf
// CbTe7=TX/9QFHP);<C5#87I<KPC+MYVg6J5/UM0+FNK:48:fWI-\WMU4RPWHT?^,
// LA?0Qd:2Q_ff;@+TVNKJ/ad:^YdUK87S=^T3Q,IDFc?AC94L4MZd&@7-&MF[f=]I
// 9a,81+&6)_gGe0@NH&c+#EAU(EEb#GXR/]NC1_(RJ>2]]_b14#^N>9114)<7#3#6
// =9OM&[W](,:2)VWfEH3Q;C>=]PXd;7:CGSPI]>V[=MTHC^VMdSA.c,V8WbWRMTH#
// ]3=_NKHgFYJP]BTGeZ:d_4b[4URE3>OW)F+KbPZO+3^2;II5cJZVdc9[[(2ITF51
// N>AUg44P<OFQgGdJ.@X&I7HF9_\6N@d&QH#Ob.d(RB;.[ZGd&AY\2[C&Z7NY3@L8
// \T+([^[d1BT-JJf)X4N.f[GW_\NJ]ZBTWEWcb5N.7)A0SVTRIAZH?#0bOE8U8-0_
// #=g,R>de6#UCVOU)@eVFX.c\aQGZ9;g_8IO?/+<.@8WJS93C-FN8@Q&2eZI40[L3
// E/?3(#.V^G@]?JZ3--ca)MQa?&7/5/CF0=CF=:Q=Q9(.=9VY+MX::QE0LcZ7Pd0g
// BeD.X(@d.O>g4,&H>9c^^.]ef6f1I[J59JTcU#Y8VZf94:OUIAS5TUVU&?<PAUSg
// .,3>0QKKQ0:+&4K5_8N^9,+3#,B:2f]:QRA_bg\DaE^<RcFV8X,(5EMb>+(#HEZ<
// D;,^>G0+DR9:/5fb(R_&_7FdIVR3^4(@1CQG+/X0-1Z\I<9E>VFB^7/^f4WH8MQ-
// 7Td>R2g<V.FHe^/F_5,;1&>G9PaR(Cge^9g8[5WVYSM,9LQ#P3b6>g(]ZJe_;4L(
// cB&E8[+3P&>5VR4MYGD0[Jc+5;\5HR8VR5b7D0=[f+8,330?LZIDDD9?1I(T4V)8
// LBdcYP9ZZ<(&(Q6C9HN)F\TDGdKX=N\&?N&(+/cD0QdDFUE6d)L27^U&ZA]g8Y4Z
// f?K<KK)cP?#d=VL_L#XccYWZR3OMCaTBW#U-3ZPM-WS^dYb(\UZQ?V:&bW?S+985
// D)I=bIQe;Q;,HdQZ:H\GUC)9a.LR;H>\V+Q=N5FcL#Nc[^c]FL:Q+[)L.SBOfL#@
// HW0A)KB>cV3[K-T+YD)&7+Hd-Z02D<+YG[<VGfAE_a&8#XNCDQUYd<6-^JAW76)H
// 31ed;6P^CPGdG\\:C^eBQG6f[/_FQgUb5g.--?W<]Q>G[#)AR-I>]B/2L[;6N;)S
// Ze^S<N2=&-9X_BR]9&N)^7QN[HJ<O=Ue1a_ZQO\Gde;XdPbc9c)TX.APXBN2AF2)
// 5E9b(85>3[56\_94@C.L_TR@&a7f5aSM-?UEg#0?7f[<_f=\=dMS^MRBXBI,b97\
// c-#Yf7M:)#W-]J4648>eJ/E)6<##<>7-DGKEaPg&G?;TS1OO@GRF#<S42AZ+..b=
// ;G4?,T1-aDB9^c:17??5FbZ(MM;C\\:BJaMdB=ZKa3Oc_:.J;Q.-X451JP+]=D6L
// 9[Ng?,B_+XO^I@+<(?]g97d>,WS[f&-CN5fe9)=5;_)UdVWaa]G7>P;L2SZcaA3)
// QS0R.[Q;c_@8ZB:<__LA?HM;2_/Z]cWS:bQ47Sg@K2YS>+7SF=IddZfQ>29bW1<>
// N:\g(.3(M?89W+4M<4VB9(YA6YV2=WEEM+/.84&/e,BJZYE_N\cZ5N6?P7>.cgPQ
// 0NHMBee)g\DRdGV.T8G[FGBNR/V@F,Z2+PS03?GF?J?dE&C222T>TA]3NO_P6B;/
// [Q9fLXCQPX@#&e-EB(f)&]R28&NB,]\FG&&]D;H]15/?eefFVH-d(;9U&</eb?^W
// ;JK.[[ZCa]g8JOI3A02+CDU@8YL\U<.I/7LKN3^-=[@QK+bX9IW>+Z1=Y3.7A.W;
// G@-UKf>N>=GZ4M=?R^c2+LOb?P2Jc9dN4fI6@bd1D^b=PKQWV2EK-)O<cf_ULf^J
// H,;U.F5LKWL;VMc,CMUK.<d_75[M-[/cg^0+4\CR]eb)=,<Z+?df9fV2-<.CZ.P4
// EB60X6KgI+b/,e6&2DD3/[0[(g66fPb\5QLP?XI56-A^bQ4NSI42A\N4U<-1_16P
// 30.X7ea69g6e4d,J0.C,>g9W-3FMA,X4e:<R>BC.ZWK-_Z1&86<SVcQ-]#-CC,KE
// (-L0D<7:\=6Y7B4ETZ<1S_O[N@AHNPJ-#/?O<:(L6RbQQ[D2_A4b4,6G79f-W4;W
// ?Y9Y=M/#HL3]Y[b\1X#?+])=ea-NS7Pac,#G@O]dC=&Fe:DcgWQST-f>,B;bW4>_
// eXSYe5CJQ9JS9U.IX4@@-JeId+[G@c;>RCd20aO\Ud^&^S^SH.R>\FYR@Y#F8JN3
// ^CNeUf>UbE@?De_S)ZF.FbPQ(NYb/YbPA#OSaRM9bL/JB9I7ZC7DLFU9TK]V1-bU
// S,?)6@Ec0:1@J&A<L9]FQC-DD>BZZdN.9-bR3\#\Kc3E-DbZIC(9-cXSRW\M]EdY
// f3M>KP.UBK\Y2D1[\&;HWO4),QS\-NW7I[b.KT,2e;^(EQ[?G:U?9Pa3AB&(ZWKR
// ]++]GdYB?9:PEO3LfL_U>Z1Z&2^I[N[&]MV2B]D1XB=PN0?JX8#e_d&EQUQ9\<dM
// 8,NeHbBWV&1KI<GC=R^[TQX_?0.cFT0VAd.W4a7^#1NR0D#^dZO>RYA].<5(-.39
// :0M@WZJI(Bd9.9^D8Xe2K:Y@M9E@eBCf&Gf@cA\3aV40L8RTG:OFU_FV@/=[bE6=
// /Ye>953Q3)[X380-aF]1.NGJXKdf]f4^Uc3=UJ;NRe(<I9@(^&BNd&V_f23Yg4I,
// R\R/9O+^2=Oc;3@-?gKXXZ;LI:eOM?ZV&ac,02Y;SEb-2M(M+&1b#WO1Z>(K4AW_
// @dW>C1HOLc8Aa06?)82^)F1M-3ZZS_@,Z(GB<F@[YOQD0fY;=.&_2SC?2DSb3K>O
// )WACL6Q44#f/PeY:52Y]_^-:CUAFJ)&,#<Q_0>L&.bU[7>[7])?#EbQUX:HU5cGG
// QIFK^H<1MXI0B,AOJ&)a)2V0TYTO,?N7>UFbdQa6FeQdINQ>/,(?H0b1T1d_>;ed
// QJH>:VJ.?Tb8^5/I04U626P?4OV-_NXP=aebFg[8,8<0@N[[T?129]A+PK\^EbOJ
// -:MH::89-VC35^P/GZ&3Z[WQc:VV^RP;/FaO30IPaFQ5c=O;3W93_GL];]E.U\]&
// 7(_C.&C[HdAKN-SH[Z6Nc:1gaO7H\HF:7KGAfKYB][U#7U&+gHZa+.,Rbb@[T1>(
// 2@?MOZ>V(aW&QBbI#>I=1)VG6:U4LPS:-Z#d^5gGg)QW.gAS^RC]5V;#MU9?LC.:
// >(9B>bW,)TOX1@7ZR^?a<:1[gBSU+.2<R5;]c9Ia,97S_J>PF]W>(NY:.gU#>Z?L
// 23P>eU&/_V#@Z#a_Cb3.LRe=M+Cg[CE84(18g986AB^F/Ce[-bKG7bZ#>U/@aS/g
// DEH0GE3WFON4C<KOL1PG_]9)XJKaD=3;)+)/-SA4D#Kg2;I89Ja.>Y@.L2?/KU7b
// D3]A7R7;H;dc6?CSM=71EZ>:a9MH5R#V9(B9&5T[WTf6N0^)1[GQVfVa&@QOP](2
// fK^@C4B#.W/>7:X\XRBB^VF/&C&7aXOTSN6J;FfE]=/HQe1G8\XHPA7&b]H82(]>
// .\M.AW257VK&QY.ZNOT09T=6U)FV_.OUbZe::+Z4f8(N:Xf9e(QRO5#63d:QKMK.
// daHD[QR3I7.2RafQ=VIg^/4eg_)9&+J5O\N3/Z\^^eOKNCSK4fd]22^CZ/J@b-;(
// ^8H_Gc3G+5(cQ;Je\HAIRRNS]4QG_4-e1P_-SL[eF+_?_eYe,<J]<a[Y3.>-7[Sb
// SP7T-502B;4H^G_Jee_5M>ONWEe^,,8\)OP.Z^FVa7N]d#F1\>)X6E#OX1J9B)[U
// :6T_+>41^/cATR-C5LeS1G6fK?.5eYMgY21_5FM/=K8)@:P&4a)&4bc0FcPI<d]P
// ILN\WH5VX,[S_<Z-e3JXHc::1N.@7CR^5BHOL17T>60<9BR+A^MHc,:g6/=K8@=M
// GHdCZE]:EeX4gUR&YQ:TK@H,BN&,MA#A8.O\,V,A[&=,641,X38U^EeccINZC.&L
// -YA\f/5bQ71X<AQ:O4G_7c.RJVZg&.XR0@3Q04+MDYA>92d_HSRP;[>/@#+]#^WT
// 9V<>C:/6Ee+dK6.TDFbN^EH(?)a^)YZg\(T@?3:OQ;6_B:a,[gfRCX@BD5[\cYR\
// L9ObbN3(W<(G,88L<1#W5URD_#8M/.7?24cZ)APH_WC&K+,HML7L]U42^(S^EKa]
// 4?aE9X^&bEF\-Ia7,J\eWb1/777c_E3QDX]9BcYHD9P?1\<AMe:>,2fXN[<IR#aK
// >RILeD3(-c<R\MWd8gDV\8(>L5,R??1DO:I6O]=K6\WLF)P)<,U8)DTSHHS#TVW+
// 6BO^81BP.G>=SS3]8Nf.T6??0b:ZDG1+)NKV@P<Vc6C9Zd(8Hf&7#WVQZZ1?Ef@&
// ?cU^(6MC#OPB=c7CPI.;T)2^HKT-QF:[9[SfYS#cICDX_5RE5>:RSK<_Z)dD0gWe
// T>#@cZTX5_#KfSeX5dg^OK=72]&HVIdJfQ?a(>MA6<d?Y.=-_EK@_M)QJQNZ\]aN
// \,I+H<HOH&WB;N6&7(<(NbR#M\_-Q^X=0>T3fPf-[_J.ST=6[@7O&-Zd6B)fKOI(
// ^b1eBU9R4PNITdW_VFZS>RTIX/[+_79ONd7BPIYW6HZ^;VM3P5bb:3\_O)D1K4N=
// X#IX/ZROP@;N3QAI>E3+]I;MY1G/OE6T9,1EH1Gc>8a8e<MPIS,2H@X2JB]gGAOY
// -Ta]E9+Z6(/Z2RObX&f1&gQ2-?\c7gX>\#f+O1d4.;8VJ)Q5d9TY.[:27[SI);V>
// K#[GHb>Y\b0M.3C1BbB-T6[=cRGM(V,T/Y5#[3KD9E24H3,>0&DM)=#dNG)aD&,=
// c7(YYA?gM;#a_)E-IGF2+[-W?9b78=+f;I@H<MF\fa+^<F(,dA7_eB;bZ86XN+OX
// [Me:V&+SW<;bP7D&M[HI1O7;>50g2F>D=/Ac.aJ;TK^RTZS;7^29MYMH5=Eg07(D
// BTcD9dR4^)ZT+ZeYfa@:>eHP@(^]JNdT1D)CK.VC<W0,CUL(M>L/Ia)3>GF2:&]F
// Mb#E,Z+Pfda)fQbL=/J=Y+ZO:e/E1GG16J<;NMUg;WG69H7Q[e65.Tc2@E@f2CX:
// 91-6Z.gS&\>.0N=.#fIH?-V7H\EN^Q5^5/BbCOC.F=Y;E7_,]DII<c_SX_2;DGT=
// 1A?BaQY8#_G6]&6XNSQeTf8[.9?/?7=L@N\f#aEa;a,)DP,^IHe8K8(L&-DA\FI.
// a^.V6P?cCJY,9aOKH>ZT;c-S@)eCKDDdGCXE]7,2Q>a/Z,Lg-:Z3fB80H/M;TC0A
// K:1Hf:T5L5,Df56,L?0R[Q[&,52MOfOM]&1Ve2[8dDFO#GBGY9:&NE8VPQWLJYJ5
// IP??B?\=4L^\b&7eO\4CaN2a\W(F-LWEPI-<9L=-FFZ>L,R?V4,f?6AM>f\9;P1d
// cNJ)5<2FV3:Y]N7:HN)[.A5b]#5Da<\YMGK8,BfLH?;6\YM17&_IX6LcD/d.QO#N
// NaA)g>JaSEGd^;eBTN)1(9d;CBbg<EDe.J.>C&[Xag)[2\K^UD]bISO--9FZND:H
// /,UfZ7W-[M@RYA2X<BGgF.DW<.;KZI>Ddf#LF[[C?8?0a\=IET?ZN:(7]5-A1<=E
// 3d+/7+C0@;K9bDK)<e2Ib/@>+<,+,7T0.2O&Bf8J4a=14S,5H[13aC2f@>f8W_]c
// R\==7>ATeeUC)^fQYKNR\@@V6g-GP>AE>[I.3(O45d4<MD?R[eSX87g5,(a<9OeW
// \+^[<I?T-a2:&6KOPR^f:O8Ca&73-X_8=fEVG))a.7-@VMc]P_I]3d?ULP9>\eX?
// >ZJVaQNR\U4Yc_JdVJ]b@2[C:+6eQ7Wg)+RQW7:).&ENVC5O?JQOJ@BaEGa:Ab&<
// e<,ZYX/2-DZM@BfHNV42MA0=7W30AVg?gK1Y7/]Ma\5]BK6Qc0f18&QW-4+;(fRX
// g&8@)K@VB/UJ(?=ET1EWUfQ]O90#bdNPgHM\,P]0_KW&[F3WUY5?.4_V4F.(FVd&
// L,?aRd(3&:FICM?CN<_PJ<6#>,#L],@#(Y8NO.:(.)bGJ;;ZRFJ/\#E2#Q2&4H4^
// 4/N8SS;8X#E)2](7-gQU;N54<EWBD:TA0>Q3c#E(P+4Ib\?.F/WecX9?(W?L_f-I
// 14cRIPO4[/;4<e=<57D;/I)/^T(]acEE]9O++<8\^EY3=M9TH&NU3DbSaQ[4Z_=7
// b_?XH^J)0e?2Q5J#6=5F0^X)),bG<0d+(9<Z1R<\O8a]f&NLW.QR#@0<5HU&aL9f
// .&Q3TQF/L8NQF]dPa[dLV_#YDHALJe8cA,]BQKVQQELfU0BB/+/@L/2?B1T46^Ie
// Z>TLXZ@QdY29ZV0CL&\<67.5e??fF:+C]^&D5ZZ84,WMJb0f[2)VSE2F1&5JO(7I
// ,W4a:@?:8f@M3I;.;Z9+B51,U.ZOL4+Y<;)/.SGWK\G+T>@OUfbE>6+5QM_B//U(
// GeN;gFZ;N=dgeR+Q)g@6(;?M6OD)5\6XZ8=Q#:8bTM-ESeGFH1WQ2_f.&g176^:I
// dG2_KHM<(K?0fe>S==d\R;^Z^bK\IUUa<9Y,:6@HGL0[1/@AKfaB-B/M#+;C,>(@
// 650IC2PH#>#HBG\/6_RbK-WIf#c7&d<ALO@->UgAcG>^[b)5/9(bM,d86Q@NbX0V
// &3&b^G(J\ZXGe(<9MWTMd25<:?IIG)(89:ZDG>ZYAW:\#R<U,N8&2AIKeXNMF@TI
// \E6E()L_Bd;]F)R3^g+-KXJ9Z@HSe@.:3,I_IP&BFe#0S9K;1LfX>;3[&<:aWDLU
// C<PP./3b;./_f.QAgI9LeKQfd@XSaYd14=/R8=_ERBW[f0BcYPYPba68CSA?=6K0
// #Nd^U(/ABB24b0\V(5Q1]=?aP<cT,VdD+#Jb[Y>d#ZafUT=LTR3RKcBcXU8dZ@e.
// Y2Qe\CcH_BUQfOaJH/(H:NEMOe8.[F/1.NS=R6+TH1EcW&=+MLgBGAHb#:JCG76S
// E_6c<1>Q8=&2?O055AWD=K07REBI4#JACJ7KVA6FFV9S,UD7.J;f-M1#ZK)/7@>f
// Z)/=@,XV[Ma_caN,Dbd>D_e.Z-<V,Sa)7])@]fTZ<XbX4TTde3DB(\C-1(X97-QE
// c[O,[>9]ETP?#KZBRe8XK2_,_(M]X0eEVQ=L/B<<E-E^eDRU0]P^1.e[FQL,+9gY
// GTZ2-C2#A2,S_0YFA/085DU5-R_b6KI/GM^/XGCY[XF5P2U(A4OFIN+DV,Sab]_>
// g.N5A)>N^;;,S<fTWHd>6c\[[2HO1-T2]JG&R:U5VEC\C?-S7)PA5BF1c]U4ZUDM
// 5F#<).4]aY]V1^aK>@=dUf:6CSJ,Ob]APbHLK2KQD@?PBM\><EAP>,9b/^_4V#Vc
// _cX?N5GY=beS.53>+,\FP2+b65QBP=866@M]VUQWL<(S2JZB54++a_2(1SWcROX5
// d#A)c>ST3U#@ad6TNcTGJ4MZ9R:0#H/OO@eF[,W,HHX+/H\7,Z]7McCaW]BSKA_U
// NE[N5H/0eK7NMgM9g3O+D:I4&a.eOZKfB4?-JG2eQC(J1.0[Y,+/=5)PJB-ed1Q,
// RAU2PS<CcM0A/Tb\JRG0CPZd1aIFZRA>;XM=/XZS>T2VX(/W8X4)&fH0b8J[ZfU0
// V+GSDfV;QNS:d@Z2@:FA7CPPca90[3g@PC:3&7I=JZe.NI=I(3_cE>9I[c/C:H&d
// DF1J[NX<M;>,#6N8P.0QGg(##YVS+0NAM1WO^J[ACF,LD]<RU>+Jb1G[_6&3JaGI
// ZL\MTH1BDURJg3b>WQ-35@d0I+OV8MIe>Y2WJgTD)MKQN4(&\@NTNY,/7c/LI]9;
// aGU5POXd<&L),dH?#^Yf,I0O[P[aEA>)VSW4LW[_d@-Md\f1LHf<LT,cT=20BgbU
// H-G<)-FB2Q/GY).,Z8f&/_e,ESUO#CB+#Y&VNOER/[F#O<,)Xd)YLL2N^)CHWM[@
// R#ZY;4,I7UR?f/YJdR&\=1)5T_@<(DL>d[-DKSC7W\_R24A<DP=CeKO)O1W+1N_U
// #dASR+g;OX/@C0)Ag&&L]H?J/,Z3IJH3THJN<fYOI&SZZI(18E1a^^J;7,c?-HE@
// QBP:WaV&ObJ#bA?A=KaMC:Q0f-MBWV)NU^ZUa[eH,Uf>3a&0A]Y4+CH#B9=0V3J_
// <;6&I#.,(@Te@;Bed#49ZU73IZ]CegWWEWQA_F(P3SO6T)OK>NJ&D#F94Rf=?T/3
// ]R+>=O]gV2(HR8-Ae]E^CKaGH8QHY<d6MfVLQRbe?<1S(_c5EXKWM.R_6TE;7A8=
// B+FKDKC,X83e&V#J?g<:\[AY8L81.Q[S#K2bK2):<89)>==_<4.[QUZ_M/J\=8E8
// QV3&RUNKgTB8G&]+.AY7(J2PC#D8LQaEO^,2OQA-,U9]fWNCR:-I);XUAQVf_)e_
// BK7;--N9ABB3aO@Y3DI7.8+e7T^.>:H4;dLMW>GNFU,I6]_V2#N+TX#HOc;:H+L?
// +_T5I^Y[O9:B[6HScCW_.HF2?_Q+PE;?C[cfSbZ4OOU=@N?)IebT(]PIZF#4@)@+
// T)BXJ.[cbI\XC(Ja9U-??H_?fRFE?EXAcRBJ[I)>BF&+9/@O#>&Q-?F<8FUfM;@>
// TP;A7?f54G(ZJ@-=&2KC]b3R5WPbIO)7,4):+HI^eKN9J]2_:d;UYGPK?P&^_@HW
// Z_:<RU)7/CI9gUQ:+N??S@?KGdBcHVQ)d^C,0/0E,b3J?VXMK36#D\.E?8+E)HXU
// 4Q136[Z&C\8QNaO<Q&adU0&1(4-Gc[7Z,gI(^\QUDLB4FEXBIQDNa&VH5=L1?Dg;
// (SF52HHFfLAU5TDTJHBL_Od=[04:>_[;<cL64+>@J^5f7K.T_b(ad+&4@_T3T:)/
// @XF5J<2G5MLG;-\VUE6M#_M.)HZ6NTCIU;P-0Gc#+TRPefTK3SV&P>gBCb.LSH>D
// KcU)J/P,W5FCU7K;E,O)49O)GVbIO5&02&JLTFG^a,QL2g88/5O0,2>C3a=fRTSQ
// DT:?[P\Q9eVFYA.]cf^,/#QQf.4<F>LH0L#U>PB,)/-0L-N]S>FI<_gK1R5<T[_T
// :Y.:\>dO6=b4dK\P>-95Tc9Pf:A?:&T1C:bNXF=4fd:=ABF\QC\-\+>3]7Ld:_ZG
// N(#0IU8]^/F&DQcKKYB,Ma5,4)<aG>2/B.<6bD/_,bF<V):RfHYUUSHd,+2Jg=K,
// K5>M?@[fTWW?B#PgWSX,aZ\)122,H^eCE4UAc#>,Yb9KZ1,b?ZD28G6f\AFF5NU<
// Y#Z<dC8C8ca9TODLP+UN]Z1IMAJD5OZNd+O9,FTPP3#UWZ9L/3Y4>EW\/)JFb6eV
// P^5g_e5BgN[?)c2a4+F>-D+)CB8YEYZQVbRYRR_7g9;&b6HYRFVdX\3@-A,]KS9+
// TI#c3:O3&R_,4,J4<(0.L-0@M7THB-BK<]M]g50N55)OTE[&88PGP^K:3>GT[S&(
// b2BCHH(<9dRea+\)d(\BB<S1VNQ/DLN:V9ac6C-+7BaS\B4-YD-1UH<R&5C+cUB]
// 05T>8:;Pg2Z>KNbBDPSLMa^18TI.C;(CZG6Mf.(W\#Z^8\PC?/baCTY[Q4&H1+,7
// X66WP6UX/:f_aFA6.9S_^+71?WF^\&J+Z.#&bL0AN4?\7B\G<Z:/]CLD_).aS3f=
// J8ZRKR+<R/N^f_>R=GQK[ORVQ6,&)aZ\E026fDf=6SbXJFK\fVD1S]?c3&M;PE7b
// #0@\eSB^[CO&T?\aV)D?F]#-\/KG57<VPf8F89V/;S11OXG5DKDb/+bA[1;RR?;0
// .f-E6VS^]DBgbMD2FYd&KAbd]=JV#]YNWDRWDIX.\G.X]?fH0;GS6=8P#717<aaA
// N/V@4L7,[@Md/?>_Ze2,e\#cVe&&J2H8A6=[e.EAI?H-cf[Z#;Q(D+OGJI>e=>C6
// +</0Id>O-g\RBY,,ZO\F5Y&ZKOG+XO7U0UU@_;:3A.8]fe1H4OOLGWL9BN:SV(V+
// P7EIaUYW5e[?R2(bERA08EE_KLR0f>?f4@0F6]-:BB_GebX/Sde>^b7G:BZ@L5=K
// He39/NC\1#[_>F7>F<e;DKZ,E,\J;Y&-?9XM1T^&.-[A<eOFDbN@+:,YDF(UPNE(
// 70M<ALg)HOHJALTI=LMRYdEJ,X\<>=?/:Vg.)@d\.G[@EA,Z1KA2F2P^ZFY\._Se
// P&^2eYUUA9CW-&BQ</=JKf7@+.2gGVaaa#0,J/_ZNaB#B\CefOf-H&Na4)&SGba8
// PKgg1OCR7a?+b)TV,G#f1JcNcN;&PT5.E(=6QU0TeHB/S)WO&7SNfQ=O+88E#_7\
// &6<+=ea:\AK0XM_6ME6T7@IE0[6a<LK7N_0:e)K8U\UJ1?RD1\3Og+?)L4C?7fNW
// T/K3;e2JS7=2VSbYe@D-RWWMFSLG0OE,Y#:bPOBVLD0MaU40I26HEb.7Y6(Dgb]P
// .Rc@51_>1b2_1XT:6>O#DS6,,G/=\JZf\cT:-;=g&P;-P.75#Q=+R,9O]A^Og/CR
// Pe26;BMF5HYI5;/d1faV,H>NRO;LLL=+6VZV;T8^KIXG<-,PV3_J@V.GX,)<^Z,W
// c<XO:#Ec^JTW\_/2g;eSC\CbS>^4a)KcMK1IHMeMeX&gCc\g9)aCVa+3VETUY?U,
// 9GW9QSc2<0=XV<a(TU)dRMfB/,bCLLPcdXB__+aG_C+-TVTNQ]EN;e:Q[^CV>U5H
// 3J(2VJ6Gab<50(54V+05B0a1QVNL,Y^9aa]I\MO6>&bQgIf6NZQED<T9Za4G#J@:
// W=II1@UAF-M8d?GAEA\N1)E2GR;J;dA)<eI,TR#>RW9[Mf.],:Q.^b>#_PJL^4V7
// LFU0A_eUWEc6Q)D8HC](?B5afHA^1Y\C2,Y^DJ3(dZY3J/4+(W10DH5>0Sg[Fg+2
// GZ<6-@&7B^B2de_/9QcYNV\RYgHNNKR79QRJ7F6B]?^@5g<(#48CN3:K^=XBFdH#
// DW.ff<Z7@L/Z-EKg0Q1QM)b..[\J,D2A&04b(SZ<N^62H[JR=^P;X0_Wc4.I^JbK
// K]MQPfC[H0;635?+.:?249V]?(56Z3/Ta]M:X84HZ/SSK,S,O?W<W>?Lg#@[gH>Q
// =JAH8/)OVF=J6Fg,DNMCK;4=TNf#Q5MN6bEg7I(QAFZP1ffW</+ZN(]?;P;H+E1Q
// E0RaUGV6I8G@50H1VVC?EQPR=.IMf_IF#\78ROOR+[O9<J;K;/^_0TFSb,6+@>2d
// ;bK@RA0ZbSe\3,BCE[Wb;I#-+.ZaF,:5PD<Q619B:6#U/<;4BTHg13F2,;QZ0JM+
// HV^(,NWW^)+.Z\YZ@6L<-bDB:NR0I:V7L.Xd:O)AD-L-f-3Q\V.8,GIIUe>1?LMS
// b]a);<7b<BDR)<^<;UC:L[c?eZ^=)&+Y1gQ&/#D3X,4S\5PY5e^H=VXI)OSC9,C<
// .#0[.=]_ZcB:;acNK,2&S@UH8MN\V?DJaGL8-3;N#=;56-ZIFgc?87+^4c3eO327
// I,1K/__OfIWbHO5::I>Ta7R1BRB5M,182@>HG)NRdX-7=VUa1W^^D\R:f)QK=)]C
// M&MJFM]<T-X[DgT#dS>,O4H[4#)IJaP5Y)6I5)-?;P77Vf#D23.bS5#42G),8>BM
// ZD?C&Z+Lb0]0/]K=^Z8#Wgg9+,d,bF?I02SY2[]ZECf\=E;D+7@B5TCJ_,O]=+fT
// cHLbFV-[\0_,XD/1,#YWW+Z,bX9ONA?IfI7CBT/E/#R):^8YJ5LTd)NgLQ)YEG0U
// Q3<>V8YbHI4L&aTPZW<?IU#_?(R&/LI-70,W5BG26a68[gM_J(Yge,OL@M2GWE2(
// R(=VR>^=AZ7R^Lf@.\&Eg2KZY:H1H_GXCdR2[+S\Z4gFS5cfCX5^e:E0Z+M5<f^>
// ,+&Ye50DcTbAIBP,@Q;QG5ZCcP5bX9ODdI2DVYS2@W=CPeK(L26#:(RKAGV8<>QC
// _5Z_<0QBgc401Qac8[(,aAMZg_+I\+D,PMS6aD8<OKCU.Y[,B#NZP6W).:^&SFUd
// @OU<S8?9?=,Sd7C^a5QU0Y6c,3f<S>HHeS3NFI]EWeMQ.OEIgQN(@U7gMIf\Qd@4
// ?JP7KSM?O<gBg]Z4GAVbXe/-K>0[_WKXZH3@F6XGXUW2.C&.?<&HHVR>R36N/Wfe
// WSYNHHCYdH=a&-BX<KJJCB9RaEa5-WKL<9K<WH54,;UA;L&VfMD5gAS:-KF--JN2
// ^S34JGGR?Z;91cBVQ.a[,?:[PI@)-LaU]EKYV;;[=.K0@1>4Z\&d33e3KHW)>5-?
// &/@e,5,Pa:8?<1G90XQA</FEFK)[H7E-CT>\N)W[/b(IPa3KKJU&d>#NBfHMf9;L
// EI(S#](2J754TG6\3AXQJdF:2]#&KY5[(2XXc7JOBcC3B<\/;_aT9QKA64bVH^bD
// dY9bL2D^H;YbIEPcUScJMD_T9K=ge9b4Uf(>W<L3?@G<XZ;\CDJ(5?I;+C\<?IC(
// ]/:WK5aR>+.;dY4Q@fQV83M?Z-U-VO__J9)&1B5+/T\1[caU9H0--(>cS[6-@d<c
// Ea5g8..:@eE]g7IEG4eT4.+11J2)U](@3GV&,Pa_JL:],:LRGZ5gDN([]RYA?BaZ
// /<50MHQ#G3KbcJeAQRJ>[&B&9c-,Ie?S>GUEf_S),>>\3F?#T:dS@2I9N,.R;S#N
// _7#Z85+;Y4e:d(2>>QQVNGBGB\EC)/4C<?W7H^>/fcc(_>A=_R78P]W\L8+Z5g)\
// J3MaHX_VD25E+WXQ5Y\LMH)0dYT)E;K#:8YORBa1?1[<HOOYg<J[;T5G;<)>83:L
// 7^<Z/[NLLM1BSag,G5[&CIKW)X9N-3gKVUPHAG4IR+g,.a00GcYUeCA3I3(?Mc+A
// <T?1e.:5[JP2efKQEXYb0<]KMbf0S1,Ee]6_F\:#+eM9R.>bHJ#.5eUe9bX.2XGB
// eE]?/B:a3gA^VaA_;dQPD54=FV<]:(gPeeP_B]8W1PB?3PZ(NegP4,;f&Ef7T]]>
// XTb6]bZY(>?cZaSSZ4M+NB56X=>Va<A_4cL;K@?S8?bK&&V/;Q1JX<FW91(I>&9a
// JMB8dOHGA-#F&QPLFU[XTD2R^&H-&KR,cd5&E8H48Tcd@H;)I,3(M1)])\IHQFa.
// ^BEJTV@G.@;_#],SGV0B+3;XMEdHcfKK>dGN++5WDRG1g(4.B@A/?g^:I)[e+g?-
// Z/?CXeTNYBCYb;,_75ST53+6CPE=e.&DA>Hb/cH^1dNaO00^5<-Oa7QL2E\K^bdR
// Z=(YJ1WM?A+;Of@X7UI[=@92F2@VCL>AD40XCgQ;^XgB+(a0+.\]R4P@^299>6<d
// OX:WPf^eg#@E8<fHW8<,[GaM#AL:?\)f:.AG\CIfZ\Q-b7FW]\dDb;B9.2BRK?I2
// ([(c_;+Y,a0:[^J;/F_?H-Nbc+H2]g8@]2,e1_K:##Dc5)UNCA@GRT2Ra9BS2TU,
// XLUa9;SY^H3(WAB+LP1(dTP,^g-HFZ^9.3,7N.9P.]G9G8ZOfHJ]9C4TT)9]WLHW
// )70;&VdPU<0;=fMb&BT<SR&gGT57QD8>A>6B8YVX2K(4eK,81gQL8DaDGBF<\6]d
// _e9@[(-HV=,V8e4/<Ud&=BUK4)^<4)PF3;?<UYeQ/GS<B,L_9,D1V_4b)8;HRSQb
// 69SE&cN&69+R#b&[W]X<^Z48FdXK1U__OSH(2Z^f0A>W[G(Sa,g_1)->YC9(3BX?
// 34F(+O7BWJ_YE,bZP/YeOf3I]g?f[O0=bH^)AaETa,D8F.XUWdRS=/7A3c&^a3)[
// K+94ZM4.=T42SRR9<\P;JZgfQXB;.QId^#NG++c^B]Y>\7PM;5]A9T>2f@bUd<H^
// 6<)[CC5bHF]EBD;e0L]bTQRXI93PDFZBCGQLJNdb(.=.5DH1G?_W.4XBI#gPP6fb
// :R95[VUK3FN[Z@:/_78?.6DC23K_^/^2:K1+LfES@=,bKF+:,CL]\gZMgeOX/T_(
// GALSa<6:2?-E+<15dIX<Q:N5M[9@FN@;#U12>DDgHO,?W7e@PM8I@V+6+DI(M2)G
// .,ZH0Vd7_M?f3L7BZV/?BLXNT4<(XO:\C0]@Q=HJH7V60A+CX1=LA0Rg,-M^8(TX
// +6\/Q9JFdSU0KLG-9AJ3+3.ge2^WEg(H05SE1a2T.8cD\THeO)0A:MP\OW6T37+P
// +9=<J6Y59.=;V.1I9]Db]\+2-0?_f]G\Q:;CSWPdJY#>Y;\5RE-=;[8gGOc5[Tc5
// >R8L=>_EYP]VU\\6-J4)=GfC3_bLF/?10#cADGWe^KSJ:>d,T6R6^#\Pc9GYNH0P
// VWd>:c=cS7Ng1,.9b>N<LL[BfUIDZ1DSS\\S]4C.O<H=?\XgK_cOYFL#Q#^82/TV
// 6=L0YVT)3OX@93,Z>)&K1(>G7aDR+6_f):U_(:LM4O&D(g?H(cH9D2TC26S_.MHX
// 1<O)QJ?Ee-#C(a/=,GT&M(^6;ME=6KR?+]UIb#dARXEJU_+)B_@NMYVYB/_M2:7T
// 9dF?;A#<US)gN6\@9/E6;g76d[MPX0N45#;9[-,127KdXI-\E,G6>c?I&AE0Q;c6
// gg.0I&1G2MH)HBc?\DYW([-SE6F]eX>TF5JFB3B3EL=9+EVM&&2:766(gC,&<>,O
// P7O5I8Ea[[R,(D&NgeDbb-I>,+MSF@7JT.C&+G+5/d9G<0fdc(3P_KH7=TAWO[BI
// 567d,0c9^5-WU-E/;7+G\aRL_:>C>:d:[F0PAW8=35b7;PWaF@WIfL_R50D&-NPI
// SK6V+Y,INaK[d2g<eTQ2G_]:XIXGP);3??YB2QbQD&#Ye5C2^B0FQT_=17_<PJF0
// 8LR]H8^fH/N\+T<a]8&I+AXSAZM08_0g(&\H^X/&L+N+M=(]/>).]J0f61B6a=.W
// KFP@FBDe-Y.>?cb\eb-VEZ_[T+9-M&6[0ae&#dPAMU7@Z9e3V?BS9aN8K<D00cNQ
// +184_6V.YHF3Y/26-74c3;A)8a.69?1b73WJ_A9++#^3=EIEF8(fVKfI.H:J?;WU
// #d2H9X/3H\dC_DT=VN[dPYb8E]Z@Yd_1)Vg-P.R)E/O+7(0D=IRDF_4Q+VL\WN,g
// Ob1aRGYcK_>2FS_OX3d940Y@^7[e/EXM5+^VU2K/S@&RaCP.ZK.U#aV.V>;P>8Ze
// :>a.Wf)d8J.EQM436/eTQLSJWHY/6Bg+BB8Vb#UcXQ^?bFP=O?,\6YDXDOFS5Y?O
// &Q6URfOf_=R4F.M&Gd.VfY[7,+3-;=^fOf1.W,F-GWDK=JL@^dg^8W@X5NY<]J>8
// e=\Vag6aZD^9IHM8>IBd]7U@H(RUR3d5@MK\IEd(MR/F2X(-Gc7c@Fa0Dd@c0#H5
// @d^BFDHAN>.Dc:DJ_+X:2Zd_0M8_\D6aG;T(WaFT-7XcFB)#B)W3De_[MfB,EOY#
// ?&[cdY&<[Z]X2gMW8[/4gUE+5fAY:F+4\YK14L88VX(>.e+X;EH2W&+\S)7;YUPV
// .>NN)78^S)4UPL,00@V\IfacD1O=@I\#F+LP[Ea&<UTb=7cX5fd:cc^OcV,]BX32
// &&LSfO>N[.,Y/cW<8N&IaP)&9[d/HJH_FO./d80(d2:.3-YB@K]1eXQJQdI9cC0I
// #2L_\<8BY4C4-3]g0#8@LB3850\_)8GT/]4X2,#DB(_BFa(<ANRF55,-fcHXJa/Z
// aXS&2TPNN)Y>\>g69e@+V9A>DFGUd+B1HeVd[g3PgLf:9c1M#9Q<HH3;]-V9gfD9
// #S4@ZY;f^G>M-ae&3U<9LHN;]Cc\\d&8X06,@TSJ].&J@8EP6UUM-[U#OO]ef:d?
// DVG8#@M8NR4[BLBPXf._KD1A.g/3-6-XL=(Jf\OKa)X@G-fXOe\41<#EG1;W@IQ^
// 2FfY7JOcS;d^S,Pe6?=6?>JVb8g2#EbfcWZ)a)Nd)/,9aZ40bM&eJF.b>T=SS]Mb
// ?7^[Pf4MN&Rd7=3d1,<?;X>,R;R1/M^gc@91YK4bO\OB0d/TFAQ=e^@W1HJKeMe9
// @SM(G\>4N4AJD45Ifa3)IXf7V>6)_14UEXOS.O&8^7g2U;+BW8<#YZT90-GW5G<b
// dHIN9.5<A9ZebX6]7FgP@PHN:]MN,_\XbV27bg-#Z-W13<&+B)7/W/S.R@fUgEPV
// CS7:W.=c3;+cg4FCQ@6U;T9DNb<0RW0/BQ-AD<GA>PFN@__+_GM;S<U:IUd\FI9O
// /5&(0L@FQLa#?YXFPWY>GJbRW\L;0;:?6b8;1+S4CSDO#^]1?BQZ/[(LBb0[KL/B
// -=(9)O7?[9SLHQMZR0\^.2Jd\C]+1DA/P(D<[4&?[N644OHZ40[IIg[dAF#DZL:L
// =<:S2;Td#.-c<5d1<O-=S(TadM#],>@)R9=cTcXC<b5fG<O72==.MY]1C3-8Q7LC
// 7_]MK)QdKH6B7#>4Ye7EAU[XGY90\b@P<L4X4PbPE>JKCB(/MC[:5UI;/abML(JX
// .b,)^8TX3]6U#DAN2Q89d978BSD3AK5D;TRC.N+<7\@NW.4B/,b6g1F-_[d#F&Uf
// V?[QVa_:)H,/&MNY6EWDd.PF5g7f)ZWK@4V\.fdNa._E_XB+;](0[4UG+&IV_+L0
// H;@<12QbHJ2L>(F4SaZdf,=BXfGgZGA5@QYB^/@XS0_>7GOgDDgFOZ9&QL^[.R)-
// ZW>/.?O,7AD.,J)AXLF5Q78;E0XRG]T]FQ)3N?6gVe.4(f>ON(27+gQ=JMFE7=+a
// ,MT\?XQ[NeJT;?ICXF26,SD;.WXT0g8L&MHH:R@BNcb.[6J8TU4IPfDX\5N/)#D6
// R6+W?#]OB3[EQS1LA>?d_g:#&UPQUXRQ[?a(/M=Z<SG<)8aP-G[5OCBAH259BHe3
// W)N)(6?T+=E5/YL&17bW=L<=aIfHCH69,TGZb=.WD\9P_N[GEY5JDgBYBb_58GbB
// H.OZ;MQbdd,/0J;W6)Ie8ACZVIN09A3&DMDAHc>3fYNZC7-O9\A>>.a32,3@ZN:N
// Q(WWI#N1_P-CW]MR,1Q8LJEBM(P9<A\W:JU+5cQZ<cNBBUa[dUH(T)]SEZ;UC=6,
// <-e;HRK#A,[Y^_N?L/=XU^c[\FP6?@KKc(U6+)-0W-7T;;(4Y7OdbGc4GDUM39DC
// WKI4X@OE&A;ZaH=eQKBNX)UD-C6U#LK/#;cIX.05HF\_Nc^P&=eT5_cFVB(AP\GL
// b[TC8^CSE8,JU0Ea9eH2?/8_URcBB./52c]Q;Ib15&)SI;]&\?1dYY6Z6>AD>FD(
// Z9C@--X&[:XTELT1e\(13DMZE3cA@[Ca)=Rf-^7_2UIJFK8_?\FLU)^:BZ3>a<.;
// W].DL31cD_?[+R]FPKL:e5>d^ADQT.5\<PD,2?#0aH8IZQG-ZG,2bJU#dBJ1GX.H
// <<^&DgCO)Ja4)d2cdIU^^9;]U>)I-44MO<B,Na^d?EU\.Jd2gM<2(g17U4L#CN:4
// Ue;2@ZB81_O@SQKBc@Y;K/_<4+-&Z014+ccM=18UDX\+RQ41<AT0(f4M8c9@/YG9
// <dY,QDMeG3ID[_8S.bM=Y@geM2W(H=dS\W\2^NUO(DJ(B8&W53NP#)DP+d>U@=H:
// GX(J=UFL7-SFI2EU]F:PV4X,KLQ:C8gO(5+gA=-f(96??I39QU[cGPTJ1--\c8R(
// 0Dfdg.aP7@.E@b-MESMLH+_C;9G65Wa=BAS^,0BCDBJ1;/QV]ScQGe/3[Gaf7YR5
// #EFD@M^bC^+A50J_V<NT5QgfWS-]==;QI\>3AMC9JALT[_23\J>gMeIId#fTb7@_
// FH/e./7^QB,PQ3TXOEF3f3=SAN3B:120&)N7FL5+gfX9+16/?.E\YEMUX-?<dUSY
// (.3YO>(&DNL48373HIG./.KKH<4H\W[1(<SK:^BdI,b9<[OFY\-U>V6fb9e+^/]D
// dLC6BM\HEe(d4)PBY,a@E3U_74QP8b]@ABSUS=Uf?\de_TJ?A/OFFF]9bHLbB@4Y
// eQA+B8^[V@\99;0;_L<Y(cdeEC9C_BDXEPcY&^)ZKa/eb7=42V28c:,CEM9.(0U#
// QY\gF:O_D5LBaWW<+,:T(/^a8PO\E;;W5ac0W\W_FM04=2,P8LOO&G>R<G8e/:(1
// )#Ja+FBO6Xa=X#VE?;ba[D;Z;VL2X:M_L0;<W@LZ_Wa_XfZ&A9e[OZc^Z7CKX?[1
// )\=UVV;(6KM.@T21\-BISI+E\6dPKK>DYCR0^+&@1.>3B20fe(:fAU8):J..YcdK
// +/\:2<&C7TC?5O@0S.g0b3g^TPWJOLI;B5Z.5g&=0GRQ(0?<R@>B,_S<W;JB=-O,
// 9GDXIc6[aS?)@YDQW^USIU?D[(2?=8d^3-CL54Q_IFRLQRH)6</CAf+WMc])We-A
// -e&3RH9YZGJ14QC_9P2)(abD:VAT<-D]_Q\DD]AZIN)=E3Y^FB?_C=;7B3)OUFeZ
// IMf>XBAZ>7DHC./\(>J904?.2O..bA.X1DMDgOBC)^@?V-TLE]&c0&_C_H(?8,Wc
// @QXV+.d8HXK^<X8II=F/7;SB@E.9#H;N],#b@HId>O(TF4eLWCJZ-NZ&,JC2C./M
// BI43S8X5-BLa.P0UO(5da6.WI8f(dL3+6eDB9WQ#g7SQ.GMEN(I]08>BLUL@b9MJ
// ^/@d&14M3(FK#dbbc/Y6T]F(EdCRUF.M>W;[^;2fa7?fd&>L45Y^7NA>>aDO2P^5
// TYG)7VZMERdgT4b^36UU&RcR_)Z7&XPJF7\NV:OS=1La@U8]J(@U8Zb/]2Ac,SR/
// 06g&_BcV3;E9VHc6<dZd.)UB>]4[_a)[-(&YQ2^4@=W,g\)4AcHbMKR0aMY>dG3F
// /c);KRY?E7L_JGg,-.cW^0G_bY[G7+HLe[K>aR]];<6f/CRRYZ[)9+aAGdG68SD4
// Q@6dEF8],^JV2XRI(/W\EaZEC?f]R-^?,4DKBPP:Q@gg5e,Y4P7b(\RXN[5UO6RG
// (6)?\Y[MSb,-6e>WG2G;.)645I7Wb)/Q1Wa?-XZZV^XKM1)EQ5<6^N5084+/dcLP
// ]0XfQWH9YO-b<_=;<?2AI)R<ZfU;L&4CdMRRQ6^(NF71Hb)4WVNVcN125K:@E1T(
// a#EAESB;D\2G:+,@f+/<CBHJ?RF1G(NPQ1IbW1U]&#M@I+f9_52/4<,Fd6Df4:E_
// E>;^7eOMN=43TX1].P<@L,D69g,&FC7eeJT=8=J?LfB=gV4Z-aRPZ;)D/B3=F30+
// S?BTc49H[U-0^6?Y-7#W^AEPbK76bJB4P04=_EM/WJ8J.1?X#1A7XTcFd=)-Ga(g
// Ad3<LgZ[=@dYI)&D:,&>X=[#LSFK(:37)I55B?eY8:d9HL&CE(./Nd5;7LY6CAZf
// bF4(&EHe4BR/<-)U#@+cO422M>AC0NETa)YT&HNB)<1GLY44A@Wc]]PT[a0D-879
// SOO)7\5-bcbdf9Cg36ea6,0b(e963N_f1+;JMIS)5M=D\T48VO(>Y4-ND:1H>_BL
// Ec)6:P+M5CQ1@5_U,WT/7\VDBFAB(-<M=A1FG7:EW6N8a<=[GO1gb8g/U?BJ[OUO
// ..1g3AZ28C(1&d6Y=#bCKP0013_3-KVHf4=\P;Y)[NBQ4O@1O/=03[1A/K-F;])N
// b7_1[AS5S+&>FfDWCBaTUbQT;3de:=R30<a0I^S2G@2//:eSfP</A&PFKeBa\[;>
// 845W-?K1^#3GXW3>NPM,fS]N1A1E^<PSc[))6(RZD\D-LfUPEI@8a9YD]\@Id>W7
// [/])bF5(A/[C-ga6e8=+0<?.2-YAHSAM@HULU\,_L1+4>7)M54.G@<V<<<JVd@=(
// ,+#V=]S[.BMQAaP#(#ZEH_V3:a.CG99B0;<I0WN8:07IN@:7-=DSB,P>Q7#R(@<Y
// ],deY7D<:>LD,C-87=O@/3Ee61I3dd4(.E^W^G&:Ib&8:aP2A]>>4+S7WG[JYW/;
// fZP++73b^Vd#U,-3?gL-YNE=_WR5@fC2AEN;UdC6JD0?:9J@U5cbJJ9M\?,Ka]L6
// a-6d8XV1XU:/Z9X<3--7e_-Sa_-Hb,+IR/:Rf1SdAFS\e9-5d0Y0#W.H:8[9ZF3Q
// PfWH>YU)CF5GG&Ib:PgA@W5\44@:VP=G=#\2M+g&_J,^:b.KCE\:]S6MZf&(1,\L
// O7<9-;G@]-@Q[D49fLXXUGaFCD[X2+g6-368a+#W,QcB;aW2P^H6/5#K/P\-K52<
// T@80<0B?UZ+1S@VLDXSfMUXL[bP.UTE+FD^;Ma9K,UCYG3J65FLE0/<Q+\N/3]X[
// Ig0ESEfYT;.FE44;L,g:BB8bcD_?Gc.>g.e>d)CTDVaEXTL]gS[_SddND2KMML)4
// &1YW2TH02-/J816YP(2e5G6+QTS9\\A\D5aL]d63?,Z\&2;^)VG)BTCVLO=0(W;,
// QS9c?JR7aT(.d>Q?V()#J8fH0]2_]QAb5T(\Je=MTB#D].210\Y=9K80IfPENV(g
// bHSH)]@&>^WOIQQcg+1,;a?89Z6b/b1@H)eAb(WF_O6=@cC/(LE4QS@YDXZ\f(&>
// 2+8eGC<&3fMZL\cd)]e:+cBMLF>8UY<4FM:GFI++1^f35RL0/4IG.2&KBW7,P>7_
// cJLgNIF&F[RUE7&MS==cd#KA<UG;,Df?Y)#cBY8)>\MBLNdf@77O+;0W;-6P&f;Q
// 6UDHO>FgJ:9)Y17Vd&-/\U<2DJ_8_+YH-ZVfBXW7K@[3-2XOI.FFKf5ID^7EA@@I
// V<X\Ff>AJ1/8E#d2LaVC?+[2JC)-0IPCAb+];CDfc55L=_+R?CT4.U^aE8\49H15
// &4ZW^:Uc;H(M>YZ84MGgPZ6g\AQ/8,4J;?-_^[W/-RHAF1@.(JO7K\\3QNF#)Q49
// 3:TMg=H9/_#-OgDJG]Z)CLX/.]XD]H.Vb]CK;C,97A0U@c\2SOJYE_f@HeH\5#3E
// DJJ(;Ke0NZ,HSR1EOH<<VF_>dS\TGBLKB#)&F[2DFLad;<(YZBJZL7-ZHa&C/:)b
// 9ZOU4KRH);9;)H5UFdg0QF328)gT0@4.\IY]a>S[35>JV0Nc7&EOMUV>]8TfO7.9
// ?4^;C0#09bfMHFCNDf_dWTA+GEKL3Z)I+U>,T6;0-+K\N?7]:#daC+-8HE;GJ^GF
// BP:(+]W+Va=LJ07&f^L39&+QXc&)OW53d/e]ggDVTDf\@,M:)Q:2O:L3HMaaEgA8
// ggg@Q/+^Pe(^7#Pc4XU5([7dAdP\A7U.&1H7\E(24e,)e@P:;-2O-=P60aFX)]#8
// 97TO&7/B^#?c&<b+OIN6f](\\2X3=.9bUQND12-2,_b+.:?f?P-Hf_Deagc?JIM?
// 0H(5=M=VBW2?g0a]56fH1TG^LZRAWUTHIBRbX7P=,47^g3:c?8P>).gO)U))MS2X
// f1aDMPF]&D\,,gb+OL/],TUI&G^&+f(Oe<&I3#[/H#/+7.71EY8<f\d:d\XP[=#X
// YQ;=Af0+@He:fN??gG?71BS5b9,\2dNfdQ0<E@L6,1D1F94VXBgIK4Z@T8,1B7NB
// MbbV;03@Q]6^a]GJFQ@d,B:ZA_bYKK&G/b^-[H3?c-U(_GSgY--GBA:\g98(:;MO
// U=#0EW.9?KHP-192,&NWP5L?ZN9]TMSXWY-g<TG5b26:YE5=ZfHTcV)F]T+aED3L
// DHR^\>>+0_)YdE2-&[<VK>g16?6d?SKDCFe4Fc/5\OJ&M#&\BFG-K1,UaQ(W4-7b
// :Uc]a,FQaRMY.b0d&dLS5=f[70.EAFKeNgF8TK,T_>PUIC<>6STe_\JSVZV+R)V\
// 97;<TNHL(bBHb,eD<(\@LA37?\IJfS<MYd1Q0EW?Re^B:-.3V-)ZV1(&g2[IO<.d
// HT7AAH@03LXM-UV8Z(YL34.D,.6-[\@DcENUV/_5+>SO]2>_A;&K<</44(Q;O^c>
// <NVT,6D,Dg3ECd]3A+LeC1(1]I(B)O=\D#[?>gKNY6SI:CZ@dV1X,4,5&V08#M&g
// :KMga4@#863??/?94E+d7VAB&TYA_7(OWCR9P_UFFY#V.(J@83MMC,I=/+148c,G
// FUIV&^DA&N(LfU+0caYNV,<c_[=HgO2R\COJQA?8>2S5<LL:RAQ&DU\C39(,0M2J
// NVa83NPX:#.-?C_T]TZOdOe.@.7C6KH\-=NDIaH1<&CMHU&:a\(f)<2#E6]KEaEM
// d<MAT.b#LSXO=<PY,=EIXUY8/[/<?&X<?RgEY[/]8dQJHY8_^[4=EdZHAN-gLcB;
// ]TI&PG=&0I7X^6:9NY<D#Ff2f\D4+^,L\:=BB5@\L3OO#\F60>1_A/3I^F6cFIP:
// S/[6BT1-^H?\=U5L)YH=McRcQ8d;^ED(&UC?,FCe/5IQ1SQFO<3VT1D(=R<C8LXU
// 2Rd\PSIW_>-&=PP.bZ#6Q#Y1+ba];Z)&2bQ,2HZ9,@PZd\]L5X#M:a,P?ONIA?)M
// D_-E;7Ge62BO@.,;4=eVg&5YcC^6>9ccW-1?W40aA@eRQ^Z:)A@,7HYeB^-+XTV2
// G?\6B8>4Q7&-[GGf;&&:VLC:Z]0e@YJZJ&+>A_@_(ZJd2P(VE9(I]85)U,6)a1I-
// -:^@7KI:F#=W.L(U-X)+(XP(3OCN6.PU6:H3f8Y\++#dS?LF#UI)0O.O;;<C&V,F
// .UVYLK7ZMVBHge\7b@60>=D2LB<FT5Q<a1H[[#8FFQXHBT2N6X5WJ8Z(_0]W,AL&
// 8>I,MZB;-X9NXP7WJWK[84d_:/1TJL7MJH^FJES<@eAY9WWNF-910<OZ^Lb]]4V1
// B:-K]Cb8VcWdaBMEX0ELTJ^S>VgeR#W:HcK4VaMa?<UJ(^aWR?1<PeK]Ta.0KP<7
// @;5PN\<-J112P@dVVL^E>&K#Wa#Sc>@NZbP814f0;e,gR&-9#:W,</JHXWP=<(@V
// 2=g[02\V7A:J8J9/G(2a)UP[WgDC+.O;[O4H8YM7UCCd1d\(11Z04W4<R03_,IV;
// 8T&E8C]Dd^\JP:ONM@;Pd3ZBUJ[.Z7S,/Y-XBWKG;Zb5H:7a,WaZ,F140;6J?)),
// FGa:87Nb75@cUY>B(6/;:D:<GPb5KGFRWObKY/4)V#<A/gG._RO8JV5;Ra.BYaOe
// 6)NV/AWJ:B[]O]]J]M8a#<TQ--74ML2-_&]DQ]Z;+2:OBS\M88R3F3]R2/P#7@7=
// A,0L]JI_]ae1RC?9_8:1He+_@@X8)8/_AWUNWZ8Mbb-I#/0GG9,c+FS0d7Z=\;bI
// 32T71)eX0L+a1f66=73[0D-457eI/S/g]X<0GL?=Q^VQ[>Y?0XbGB(?/05,Bb)[A
// 75,:/,WLC6#RKS9<7KMPWBIRb#EcCDK+]+cG+2AH[+UaTd>?JYg\cX8M[^IeV3IC
// =6KX,d7:DU(2=T@5BVB^e83+-Z/CA=4RDW;[1(,Z@QV<T/WT2::7J3;>I>gd(gLL
// &)8H92CF;F3,DDJ,EgY]T;EfKH#[=M=(S,.OYdV6C]5Bg.41)X+MENQ?;:Q6@5Ve
// W3GQ=>#THIIBa46Z:+2JM#d[40f]XB,2#7-81SW4P-ANOM@?#;A#g>F<2>AB+=,\
// ,RJ\H<S8U;OLI(1:K</g,I74;_e4)HC;AD@N#1YXN?9bc@B>3C[+98DBKJa3IG8>
// b.=(J,=dMCMAZYTKG+2BR?JE<SPfIb]\O5QI42L->EgU:YX@d^\&.&(ZA[Y@ZV[G
// 8GME+4#OI8RDB1+_J;.\fMOXf/&&+6VL&F[&:R:7.&#=L\M7.Z/6.W)]PgO-#;d1
// 8c+7g^=@I2ZL8)MR.C?1;6)00JZ6HD^VTJDLUBPKT]@=[R.0T&<4UcGHc=bD].]B
// -b\O1,I]>?BcAM8K2YEV8Q^B34;VV9>:;7I/RLEXBRMMRI_7]0d<Ee;6?De7J&_?
// ;<OV1B5RcgA9/75=A.&Q=RB_J)=OZ@T@EA,1/<CK7?Kbd+c\^SbY.7Y7]E:Q76,K
// Rg1X7CY]IQBJ+(:e4HR@N.GS_WcG-5(^]DY+H_-eO475=<bM,SD=@]LO@K?1GJ4;
// DHK-JfL71S3>V,\.HGTIe]SSG,J<S;BEGT+Q6WKL=NF.a:T=bN.GeK(U]5V-&W;/
// NPPV^XBC>Xf<FCCX.X3Q)OJ;DPFK\-:PWR59Q/E0OBQ&F:faEL?FTcV2FdgZ5^PZ
// >22EFJQZ,f_KZ-U3d=Af9gaTc5ga/@[3aRA_W[:3bQ3QI?HabN9K-RM/5W]<[W+g
// )@M9:>J=\aFE@4)<PQd_@92dJRW72E/UA-7gEAX]G\_.DIb=d3LRU<7(8>bNS>fV
// )/3N&;GKcFCP,GBbd(^<1WeS[K72>N48E\B:&B/H2f)::PPg(C\&N:&Q+b(\CX8\
// 5b\ZWbZYYf9g0ED0MR6.2KW/9XHbd0f-K\E\.HP=b6VDFf\GQ1MJHD^Tb2I]^1fS
// [YJaL2bT[9FDGDARXY:CZSY8;,D\2[_8G1WX@8LI968?Vg[&=[c07\AfHHJN8dP;
// XA<1I89FF&A^(LJ=[DY>BgZ8b]UA/&?PW)5[DQ@DJD;_CQI)aF(T;\1>:KSR^4LJ
// >M=c?8:f^+?T]DG@B&-B4fc>7)GH34A1M@8C]7.YL2P,W=W9?\=HH+1F6gVcFMHa
// gKg77IeS_S+[]K/X:O[Ea9e?T;>G3F/QEdg]=Q9NdDYf([c8[;B@D^S_P>Y/Z&#I
// .LG3(_4cAID=W2bT4Y^YD+4>;;bC;IMZVP,,,XGe3]2=e2\bQYZ3b:KCS&K;:[AA
// O9F-fP36@1JIYB+9ZNBJKE9)DG&>dN9IObU#fHbPGT4dTUI<7YITG9BG.RBDBMKE
// _Z8^_WKD-D7HLf#AJ2JQg&-ZMJ,:UO(4)^)^f>HB=6S9F<Y14?BM\A^a?HeOAM>I
// LX7LQ/3APNcL3e<5GeKLcgEHS7G6:L,NYV#VVf7<eT(cS28@=2>U6N1:L3BW.dcD
// <R/D:SgI36T+,T(;EFF8eFfOb^_5+Q#96..8Od7<DAacbYYFV90FC7X<<c/4HNeZ
// D((&:U.85QK^/?>AFge@NK@^#1H2\ZLf,/>DLFde<>GfW#Q5FD3fD)eL?_^d5=&L
// &^N&)]Ef.SO3gF>SQ8A-^1;92b:P=,7T9L+J@2C]L:@(^G256a86f[XE7Y7[^#@5
// e;XJfSPeMS@ES;:Y@SH41f]#Y6]V+CC:6g,K-I603G64NH_:,4@=P+O&<#fC4AO+
// &UReUA3)8Z/0?A^4>:B0gga/&L70gU]DK@F&,N_:6-9;HA:[5Jfe5DYW<7Vebb:\
// [YD(^]fD4]DYF@]4&c9I]::]O-?eU)?PF)R:+E=WcH>N]c8Z\,]CcY<9J;^D0[[F
// K93FeKY5WR\P&C>Ta6\3JF&US]Y;B^)3c#BS#_[>e(C:ec]MA.L,2/Z,5^Ec0WWH
// 40-eI8,g<d3YYG+VNIX)SI]A4.[EV98@^IKOgMH&&6+/U,6OZ-_)\)US4T(KRP_6
// Vc[;Mf>KRfA94BN#6P25g7>-;Z>1=@Z0#1+;f2,QT,MYO4aV5Ac&UDJcJM@&GZ<)
// T1-N;R4R&W<:/aQ=M;f:T.NJUQR4N8QL;UPN&bMC??#;?5QN#R5BG3F@.U_)KfgR
// RL_4>E4RPBI?P@T,]=VXcF1<@DWCYLJO_OR@NgCPQ</>DFfLV-RYI2]SdRWf^Lc[
// F(DZ<XJ5ZgQ2,.0e9bW=8@ZZ)@+Vg0a.5BQ/gY3X=>I?5-/HMK7_O]/D?6#:F=Yc
// ,V_X2d^a&f)LWD#/V5JZCfC00JL;TD/X>S.?cG1,#f[6BN=SX0cgH=)G9YM2EJM)
// WDV#ER1OT+KPB(e>/M]M?N(\\8/7.@Q7RR;>RX0(03b@:+XV#_ZUK3,./8RDH;C>
// U0VNP]Xg&8U2QO>+73,X5NaR.,^LYQH_cW,AY;?[Cf-]XMCQ\0:Q@RG28/=5@;eY
// :1bHZYg)RV&^=OGJ?&VMM7S6C,SG&>50J1XU#T3^U?<Eg5.G@SVa<[.aW_.f:A^5
// ?9=@ffMC_?LcHgV-UY9ZePJ><D+E\E#P3d0\E)4I90B157(37KM^J4ggN=5ZeYf7
// B,&Ye&FT2DgS?5A\5ID7CT_>]&G59Cb/eg:[[L1#fQ#YFfU<]&XNJQ_b?F[45eg?
// &9(OMVE1gd-GU6R8DYT6EMSb7.);5@<4_((<96N3J@Y8FNM^+:^YIR@S#-6FR)>X
// JORH_3IYbd:[H/?H+4&#UPQL7&\OEBQJ;-T61XI4IbZ2/2^#Z/H_+-1[[[C+C9&(
// #31?f9D,\/-<)[;?(H4SP/B=]8[]-f5_VIKJ:<0O?<W;?Yf8UQNe^RX&4SgIa1L[
// KKB2A14d2S4FYXQBWLMgBSf7[^a_/2:W&^CP@\)AXcc,)7E#)-FF^C;^b?0;cR15
// ISF/=^C6=P)P+P20:YgJ4XEZMg[b[J2RW0Fe\:[#<2g4:g]A8\0X;aP:U[]BNR-G
// -I5S&B:5D,KVTSQgJ8e>:4I6T1]&SC+bWbJ\I0a#2.L77FT62>7=(5[JcI<F?991
// c\:b63BA=?(5[81,,AUJ3d>9M5O)UMNcKUAT]XE0[PKK5.^K7XY^C30a>NQ(&;FF
// 0U/4cd@W&>[^RMTWJ5]R6N]P+e041H3,UV3<1&#_I)^-\\bE8H4YJKdG?BcA7;,e
// cSH@=OQ&\WIX3c]GHd=:62P9\.-XIJRUGbA+7TH7XT[CD24Ke9]-;HZ5=[<eM<F:
// =_P_YIZ?Y6d-];5MW9P.J^I83L.,7RC1J(&aX2<+1WB\G7IJP;/1+R),Xf.BPZPc
// 1EY4V7?2#:>4=B@bSc8P(cH0;)e)<LNC0HTO8#]9E4S+9+)+Z=Rg5(^G;P[/+1D0
// a6\M>.V_a)B&WXa;879N5URg1:OFcF=39Qf[/ZRPX3^W,(--YDW?>)\7MKK5BKR7
// =45V<=Fg.Kd2IDD4>3?F7EbM0:_?+fKT<R27-/aEZLWd^P&BC+>JSI^\0=?Z60&G
// \__Fb/#IM=2RTI?NbeX@35:676+V.8-TVPBYH4Te_AN.FPFF]0669JN\SVEGKfB?
// V+e6Fg)NU:Q2aCQ,)GW0S^GW?(DcL<0S=9N3c9OeHd1L35b^g7gL>>_H>B1O);[#
// =8C::@ESVYdLa@94YT\LJgJ@)\J89KGM2J1+3-B63D2A;OI7;fU6#cWgHHgf[&08
// Z^gO^Wd=.:I;;KWECVK_-1C,/TRU,FbS9<Z.3TB3JeV10QCge[E_^(c)4AX#]:YZ
// IP]f9\5,XB,(3F7f019=-?3:8(c.HO=](@/2[A-#2UO()fY:/P;IRJQJE<1;,:RV
// Pe2<)BOD7<Z(-E4GJcKE[7B38=0HHYSfN,;23YYAGMf9_9gYg6#YMPTbVMW3_VV1
// ?:d?+?a\Og55LC5\Xg>3SIVSbL[BQ/06/\TT@.Db[E^;8[UO.+PNN(OCV\1gg0Y\
// C7H6RZ?++G.g?1(DY)NO<d.;:&2QdU:R]57cHGeXLgB]gcEEXSWAE8YXL3Z2U+C,
// =/S3A;X01H(H<,J_L=8&,:8M+(a1&2_<BDC&SV837GC3E^3C<.P9g/a,U\G.-Zb9
// H<^8Re)_B70V7b?=E_b<^2X/ed-J^26/fQF4EM#2c-BM-U&cM>[QF;=(eHPJ#RdW
// =F1RTCSN,=\;ST^6O0^>83TO:)3F7d^T:RN.B=P17OKbTDRfRWO]B(_BgEb_f,WO
// /3G5:W:5RKe+F>e/Le<HK6YQQR70B:d#N=&_)JG^OcI3N2_1&@/HJY:+8b9_S>ID
// Z+.2&c-HJBXBH<]8/c9H1QIIDP:4&JDZS;/MQE>P,WJ>U1SQ,(Z\M.7S(bN/GK/0
// Z;&1A]U1C.1G>Ed3YF0-a#F^<:Z1>,H(O9GHGFOAcY4-7cS7TZ2eK=DaX:)0/3T(
// ,)Hf2RVGV\)e,(2[eQ(3SL^91F)9JI.?8.?17XP0JGfL>PN6Y_Q7+5+/MM;S_2Tb
// U]W/JZUSGNC=e[.NH7RWCJF##,7JF]=NcGeXN#2QBbP]FZE/3:NDXNN7e-Vd@#fa
// X@[FdQ:_=dKXgeE+CM,V\E0K=\6F?d4,Y[9]>J5?DWK5E)ER39TdV\XZ,([6XV2e
// NNeR<9HPM(=9R)X2EX-b62Q&=VTEAJH.?\V?ID,QON(N_26YTC(/f:+R<BUI=Z=g
// >dc@Fb/fEP<gBFb().aMgT&/be>Z9K6+F._bg_,:,S#OaMH1R4Ba-U#9Gfc&J7M3
// X>_(@V+QXKe9ZY.IM?_BIFO2bEU66?H)K+O5c+NMW(U728RY#R5DHI5<7W?VWT^;
// ]N1TOD;,/b1Q;fBRF+20acZ#D9]@@F+d;Q4.QBX<=c#O3JQ4a,5G8QR4JWU]&EY9
// .]Q(FgCKB=ICL36g2+UPTO:]XdO5I.6[@W4g,W66SIDc(ZE+RUW??\9MAf4I\88_
// ,43HAH4+=#IG.93MHg^G-@f@_c84NZ-9=O]<1-B,MD@d=#Q73;ZEP^J[aSMUN8]Q
// 5OgUJ]&&/g2b^B6)/0bL=/1H\C&YVE^ca\X9MgaAJad4@?B#PNH[B11bILK#H^MS
// XV=WUHJ-f=f),U_T7e0f(E_:\1H/GUS<RGWB-8D2KUY85bTQ+C:3:26g4H>FHE;7
// FV_3:>7=Sc,R6O&3X#QK_UeJAa)NB\FePPAL&0#7K?U)KG?_:G[g1IK10I+>H&4c
// Oa4N6SS[_Yc<RX^>@;#.[E?4/&-^YWSHdT[0T8.-Ag(#0U5VMeX2SIAcV,UD3L[b
// /:&Je<5>L[R2YS^6Uc;+,7R(V,@DU\.(X-8cM6aOABD0AX,P79+_/=_NNRG0&958
// Ad1e96#/7)CWf,/U+;>/d7EAG34dA[]?N4-ZLWdR\6JYGUK,U>^b-+bT<VZedARG
// N-@K\MFH]+;:X=gg#LL&^8Ca@Y5dAa_9Zc9O^DUCC4,L@fVTKYLd-cVKIV&F(LIL
// AH1H--F8P8#FDgI0.=AN_ZHeZbG):\5_\IM\c^/Bg;;f/E[ZcQD;^(S3R^^]3#<N
// 8<\VB#Z9bZWJ3CN04Y11e(1R]B)\PQ(CH+b5J#;+R67B]fc(ZELB_L,2dF2]&4Y&
// ._:Z]RZ=B#M&RIEa1)ZX/c]PPQBV\<HP58g(VZ6E)@D5;d[K1PU-B2>N_FI2H?C=
// LL369OH7-PRB)_bJSB(c;:\fa-JSGBg^G[6@CUS\Pc7NX(HW?3CK\b7(&YeFZ&+f
// B(eN>F,&6.X#-PIfgLb022O4V7D&>a8DffF-[adfN@dLgS6X-<6)8D]#5cL<Tb_7
// &b1dW3aS^NdG?NQbIL[HGRK_0,b-gGB/_/=VF6D2ZIXa\B_g1ND8MSLZFS>?;bSP
// ZZ;a:+DW>(SP:RcV?VX]dJBXWL>>-4-\[5,0)<EE,^Q5G@PLMI1R?S&BM9(@EEO)
// -Jd\>g.1b0Bc4BD<7K^;P&(]+,Dc+NNeSUQ/,2\T.X>3(C;:EM+d#\L>6(P&5F;a
// G@6@6+MML]SH-^\URg,e5FO.;C2dREVA-MZ,bS:68B:K0+SW)^WC;URKIe6=:-7<
// 84PD^\Cde@]eAPdKZ>?6@CgR5TM3+H&:c/)b>(:[gW1:-1M_R7/+e5,=Z)L;6()b
// HB^J6]6&YW]0>/CDTBZEM+Sb9P;34JRbgVN4d4cJ#aJ8]F\2;59X^+^Z,PTbK&C1
// <V723&@Gc#f\W]_C54IggBHJO7fB36FS>-@PEJ_K[3VQf4-K:MM7/>1B93TQJg=E
// ;ULUg>ZB4WHZ0+I51WeIR-fLfF]/a?62&YS6g5U]]?OEc635@P6Y:[QC\^>\?./4
// BR7#,cIHU<87VR^U>JN5:W8W+[]\H<O,[-+1Y.aX_O7:IJf=G(DM<7a6?7XcT]Z+
// 2AI5bU&CGaG\<^>C^8B>4?I:W.ZX&<6V)e2M/M?T266e^J&6_TNfZQA+,/=-cP2E
// [./<2Oe@BM/59.0RAZF[G?Z9b],ZU5P5a+-<:I(Y]\G[GIKT5(/XRYd&?8Vg7PQF
// =X.]aO27^)g>^;gDZ9AM#Z,?GfdYF3WcdB]:D\N<D[?QI&8c^;Z3DRHQX<@OMO[7
// @9#c64+EU8:Q_/P74GN]QP+L:?[V\L)\?OeFV\^IZ/;V?H/2+MI_WQTI:OI99cbe
// 5A>@?RR+Qd.-=ZQTc6:>eR33@e=S7Oae@;S:?[F5DMVZ8Q\HY367Z=Q3Y2@e^SRA
// Ug<II<R=Pf\P]:&71;>]?2BfWU5+e5JX)cJG8LV>@W?0=^=LT)[Tb.@@;=0_LdOI
// ?c3b2HV4\<@]:A4,;#OXZ@F&)Fbb57BF0.B-E47ebc842bGR3aI8)&?WOG-P4CO#
// ]GfIa7M]fVAXM^#0Tb[HQ?6(acGD3aN57P/^+<+,)LQd44,RAG7+G]Y)=AVU_YMN
// UbMAYD&&+OcR@=)UO0G9FIeA#NB4Z-FA5;Kc5/]_[bcCRJN[W7YCgHIS^AN2<4W:
// Z_Y02Z,EV]f?J0,B1=VBJED.Z3Qa<\Ve;A^4FD+@^<\C6;,SH#SgW1]HAJ7^]_gT
// :@\KU7+.g2@^HF/LZLbZ1fL>,fF@@FFQ_7=(IW3Ze\4/SMQ?:Q_IO_[dCd.[50K_
// )9bgIP+3a#4Z>S0&QG;UK?4010<@6R9^E=f9^d]Gca1=eJZgedR.=TU?@9]@>U8C
// D3?0M?)cag^C&Sc^1J58@7SV\@;Be<-1M#(bQ_:VLb:f##6Y-2;A5-38_(UX0J\0
// 5^/6aTG/9aK6E@IRJg1L5389d93KO@/B8&77J25fWL5U(T7/BV=+^.M?RA\[V1Da
// bQ,&QPIaaBN,2#TCaS15<e:e>2TO0@bG:19VZeA.g0g^134DDN@/6fIV9\e2.8E-
// TN_7B^eIV<d6D3[4.:^M(fF&X]:AZVgFN1>\<Z[?a1K/1T=W?B&&:C]4>85<g318
// +H@NDTVZ]:aODV:CXNfbN;aF8T,96eMJ\[+,>8SW6&USb@g[-f.&SHW(@273a]B<
// 1W@=?a3Y++VbR5S,f]GS3#(>e,&5S<UA<K5YQ_Xa=8OHg].-]RDe7TB>b])cbMO8
// MF0=Sa?)(,5W^^-\)P6N1FE=/?W(8ZR+WRbcd=)S,7D>.;(7.;9P\I-AID][=d9[
// 4(P&W3._Q<.B]4gT8KQIc/Ud5?=JbDJ-+XF1bD0T].7W:/Eg8\,WSUWE5HW^#J=7
// g([.HC0=E#:@E<S&^=83W<cY(fa:#H9eRZ&BO&S:ZB04.D.4LMF<e;B3+,GE9UfB
// C),cf@]aWgHZ-5H@2E#E]>6B/1W+F\I/D5df^5H;UX#^GJT?TX1D(,]N?@SBD9CJ
// Ifg_^<?0\?U>2FXW)T4LT1H0@P@Jd/>=;7Nc:_ac9)g6CIMC?g;B4)NAg@HE3B.?
// V=&^c^e+#>I2LR#J#W-XPa^^<]+^8><be]bWO89<U>GK3TEF/c^(6;9g=S9BP]JG
// );NVHD:47<,(&+QYe[(Oc^IKMc?MJ-aC>1C\[@(A5ac9>C.1&MRNJ6D/Ob/L43bd
// K6DBD&c>27:Z0_C0DRbDMAKY6aO:Y)cdbUNVE)a8#FZa3^7>&I@<B&.XE-KJL3[^
// GYX<,\SB8E>UedR(1<+/gZ\)JWVG.O3OO#7Bg,76+Ic)O.T8&:L7dAFGEH9H&AVZ
// .RCb/>bQ;0]6cQ65ZS?XSf(NG=E&U0c&e&IbOCWONeAHIUQ9C#<NRcMa8&-3;;QR
// Oa[ec)0J2ZR7RWSX0.+]:,GX/K6dL3C2JN@PC>adI\[3GHb9KC+0^3A\AdV<AS:>
// ,^CU]LZS&[^^T]RgQ)Z6a^TY.DBV.[(UeAMZ-aB5A6^T^UYM9S;6@WHVfMJC(gSL
// \::CJ=_9C)\(/9#3-YN0GeK;bZTG3eCcF&51<&FLWD(LNWV@Q@A8egace]3RP&g2
// Y@NcXaD5[c/<Yd01;WB(DL-VKaKd(H-[PZGUH?&F(-X>e34&f2&MM75JYN))QG49
// eZ?Ve:4UAd4><8_0:[g1Bb&Z,&dDH[dGd-IZIX9:YaS#B4K-])]YG,>E9:L\UP7Z
// Q>GDCTE[09\=U4JSFX746;QFSb?eU5>:TM1@:67L2DBaO-Z40.dLN^&;Y,WK;AaK
// [LUY9:HYNbB#XUMWM8P6YBV65XXICdI-C?ZZ]]PbL]bD9U5?1[.P4,7S:QBG>^E9
// K,^Pb-)MFd6Y)9IYK&.D@=;H0g=\GN.YXcg8\Q86N4A5KIHD(4@8&+fVTYEd19;S
// KL.][>/&@2]PV8?+?f^3_24VZabKP@fGO3A?O=bY<6e#^@>PF^1VN/SY]QK&_5g5
// 9-LSRU8=#bIGfd<]cJ@<E\6R[R7Gb8#KY6@^?XNCXS&RP=/QAc2&<B#(dB<9DM)(
// 8IRTc;FQO?_M?Xa(&Va1Uc@DGP_<N__Q7#ba[Ua>[U(+F^9AT-:]a.).//@4N?]/
// 4-K.J##GDe@6,3^VL(K3aR<>5dEAV#3MCMC[bEE-&33VT][gcPD=+GUUJc9=7FNT
// eCEN9+0>H(.b2fNbd>V64<8FgfIdK[V)<493f\_e<BA_:=]R\9caZ8:VXSX9>A61
// OUN7\Dcf59@E\@W39/N]_>d@Y\d:46(XKCVRE=;0O:+V39X00?-1a(84)RY=FA[Q
// A;MA(/H9/DbJBA5XW&:d]9(LK^10UMe6XaV>XO17;YZ<+&.MB6N^_P:#SNEBbX/1
// @FQ)HS_+.=:\FQ^1N-#DN70(Z]CLa2@dB+5#7(;AG6OT8ER#^]B#[=/c\HCL45]#
// D);YA#(8C,0c]+]Oa\[G_Y=5.6fLR44U2KbTD&:9F-[[MKX#I[a,0cXg(JFH?P27
// =c&2;[E?RcgNaJU]URa1\X9VW01Y(PNTBJ&Ndf0Y-[QJ9N/DX5)cU-Y3D]?XgN+a
// MTXeCdE&b/=V5\McfWE0e(:?LWQb/A26/Sc<4YaY,/5@YaYH07N9_C[#2F>PHg;K
// F+49_?G?FOAeV8,6V[ZOfXO4CFFTU^??-EA66D2d:;@A?@^^1HL-?\\VE(Le[Bb,
// ZOTF)-?c\QB#BTJ.PKK^#E&U3RXL7bTW?B6#Q+bZI.-cW9/bV#G,OFReCMQ?I:G>
// fE@@SS3/JI^c]P3\#9H4P-FX7CU(dE>IXF,.D92=)7.H9TFN\)f^5fCEc>VNONYH
// K0A0SB&O-agc:0fL;L,D2;_2f.<7XGOeT+Wb#-]-@/3E^3e.[3CKPA\@2;[1VA?A
// AH#.^_fR><UCC#_2G3[D_8ZZ>CZQEEHN\1(3B.63eXV?^_T2bRD?-:d9bXRK:RBV
// S_<HG-QUU-Aa?=adV^\0.d;K-]Pb:.7\NVO+3YIUJTW^1Z.YO43Dd(B@(C:fPg.a
// TH47cd7PR2@_/?(.N&&D8TPPPa@_>?/]AB[>-NYEB7E@-O68cMYAAG9beGeQZGXG
// IA;gSZf,c:LR[\Vb&_+(;4c<43\>K.bH<41UHVfc[H,SANVgG.U.77EP-2cB6?f]
// ?X0)HV,RT&/KNC22E26<]_^0OT(X1;^?7<4;-d?,EC3C+.#N/5N730.\[ON:=7FN
// O]M,XHH01@OZ&O-Z&ef:YdXAJ94M^JJa2b.;9f0Z7I@EQ@R^7EFM@4\B3[Ub8O_?
// WE9N8NDDR,9Z1gUVSUU/Af[\T++<T_^FCOOYUcRF9:ZYV0<4V9DG+0S.fFcWQ#Y7
// >5deRH:g(:;eKD=1ME,[E#H2]?@,PTZR(6KIdI7<5^=;E6,(BfVaYF#YQgQA#S=N
// F1TC5HFVWP35-U98-Q)#92\9[FBP4H17\e,OWE,^;X2J@&XJZ?@BVD5f:g#&U2>J
// ,G6/O)6:_S]>1WPe0VVLV,geA0bP/cSBUT0\Pc:)>2Td<F7Nf=C>eA6BeBeX]Y?f
// a@8NJ?Bb^4E221K]X._7gdPJ;=GdQAdP5f+ZW#@bPX7d]MX?&A]JHD8#C<e&/9Wg
// &<_&/f<<OdMHDUZ:U)YVJaGR+(?#\UeH)(BES>V0]9DGMVBc[QO.6MKYU=f7]R=+
// 8=YIRU,gcd_92&IRM=Yb\a5dX+S0A545I225VV]N-NRX5@-,TR5/XdIS,HX8GX.L
// ;&,V)QA-b#9DGM<?J\H0b3#S-W1c9@6JfS4f_cN@0GA^.KMDfgCXPS;FJ+Q>8QV@
// (=]JWDJPIPLN5RdLA0)gC2M03b/AE]Q.C^B^WL27A,9-T/[aLK9B]\57G3F4aD_K
// P7DXW3+\QY:-DUg^cab;7[:(Y1P(a>ed4:HP@aUZN1,ge]RCN8IV-UHD3,WU(6AN
// gT#.9T)&^4AfT0U5NH:a5eD(]^4).Sf\W,.F,G]5@9,M[XXd[,8GAF9VPY?;7KQ)
// ,<H8@TKGP_2-eXE=gL,NFY<LUd1/8b6[W6@E4YFC28,UN&O[)+<<AEECd3U3<f#H
// [4P\\WZDe]NKR.1P#<YQ@S+\FFaT<;^V+;d&5Q?7OHS;8\R1WOBPR=/Re_H<D?7D
// ARK?#==#9f/a5>J#K>#^FIVPP67WP_WMeZ3-\RPA2FB#&H73)Y@ZSSEVS)?7_4)A
// ?NYB/&611G+2&fMC_H4\IT;K.#effY[T8QTBF)LaE]OK.0<(]HHde0.JS>g(>HL;
// Oc_]J#:TH40>P-KOcA)&7W:,JeHZB:8@]9d=#]E([Y>AdW@;gQeHE:<W;PR^+5=S
// :7dB66P2+4[Q_2e<H;HdM_TK425Y3=5H2+cPH?\(U6C/_fD_?&9)NP[#?38V>eCB
// &N4aF4b2<MEZFTSc7BJ]7#_#]F#_X-(W>]<FYfC<O^=eFE#(ePfW#;X^4RbIIHK_
// P:VUKK>f9aVcJ=(,LLF311+NEUWNGeJTVII803UQP/^R<bL^1^VHJ[PH1O&WPg9;
// @59@EPd\Bd01A-Q^MWg8/V&[gY.9]K_C(X,0#2g?G-f/a2Id[^?<K8E,L_OKH\OB
// 9>=4BJMFIf\M+TKD9@]g1?_7]-D<A(>=7^Eb2ge.g91O6MI,GdWKL4?[C2738M.9
// MXZ^JgR\KGc;+G8MN@>3U(@AH2R?41g>@OAM=EXWX&@;;@Pc7\+/L56S2B+QPeOA
// [-#04Ua-Xg02S\__&eIXT?1F<5Q@>WI4>SF[_VY+c@Ld,bFGg^C4VBc@3E,Ra05P
// H@gbfS9(1P6<fB4W,9;IYVT8.KQGN7/e-DT(g;H>eWE-a#0C:)6ZbGR1K.4NGG1A
// J4-abB(=E]@.PVI?&/adEETU\=];IKJ,0FYdgb/4BJ?aBGUa:(@;Zfb9DVANCEXX
// S0L02)\F&J=Z/H#BP=[MD_BeQB8fgM_YL7F=bWf<[^5ZZHUPP+9KQ@O0.8fU[T\S
// CfU8P[6CP252?efg_J;.FK^T2R5W?.Y+=<8^D(6,L[Y<S7>7:X,TAKN5OLg1Y=\f
// 9U0TB2D[a,]3\[=^]gY(E;?6.=:f2@2LL?ZCUd;&2CB3>[AL>H[(d&a3@(gbAYWT
// @?gfJQI/=5TE^&IR:g9;gC4Ve[MT2LHa<@#EG=IL,..RL,4;OF:#WK#\QAZ^4;/P
// dYE9]a48/FLA/TYW07g^)J8bIGAddPDR0\R[]2-d)?(L<(M(>T1C[4,G9K]aY&#Q
// ?Db64[MP5C_LWYC03F/Y#Le^G\>CSaTfM#:_>gW^&U-gCFJV6@&8E01dC<\V0Y2S
// \/G?I0#f&:_a<T\E_13c]I+6:VUP:);==gH-?RcP+/1F(HcO<W?F,=_a9(GdGZ]S
// DNbB__G_b==e1_=AGaeSJZN3(@gB)+<)IPV\/?B^0\L_VY9GF-L?+ACX_19R#3PA
// =OY>^,-,0C01<F+.[N3Z:O>M7P3X/5,&M1&+FES)YEYcL=dGI\2eF[J?NAA+gV,&
// <aZ,_O1SX3:MLdd:E=HC2+7c-?0>H^YY,):\M1ad9IeDA60#N6+;>/ESOM&+SF16
// 4^DRDJB)+0Y\(P3>M[0XK/6Z<R#;]\.O43-,/VcTf5XKg[V5S<EHHS5TE[8T-L(R
// X?U<gW1]+.<,aa#f;=JTC\YI4EKa9.Z@X4=)LU:=0E;WFKa.&9QJH>P#7EX2-X,3
// UKL^f_\a0P(Q]J6<A:YZJ@ceA+Y,5E^9a7ME2Zc7;c+X8VI];AC(91Ze2XP3EAVJ
// Wd;A0^\.3Zd2YJ/D.f>/&c?)#O07BaI2\0eU)0,G?N>aEI4(Md,;3O=HV@94OT\A
// .+2A]0H8IWC2SX/>[T-6)).]:L,W(\,.&S+#WLcf_E./5eRg2SZ-W[&=XLK;11JV
// AMJ2aGF_Y8?30SgI]^(8]++LCg\QT&3A8BZOH2^52[TGdM)/6fT^>A2H0I>Z_1-@
// SM8E+0UHV405+0;..Z09c.b@5f:g-V?DGd&0@,FZ2\&4NTN&CYOYSXDXSDVS.=WW
// _<82G@P34\77NL.:[g2RH;1@W;S1ScKH@]2T_<KS5JQf1V;)43_g,>J^71]1.Q1=
// R[I.dfc5QfXJ-f0S<FW3P<Ua+Ua7F3<M\,+?BDfJA_PaG[PZ?/fRF/QX]Kdg,6OE
// (@5gC=)W\dL6^g=))(8QNa#3D4OTZTBK]IOC@fd+)TAZU1E&:Iabc#.\aO7^^JD7
// IH7;CaN8>+CXE9Rf]a\VQ+N<52I0H4W8?O[fH?5=\_ZE]/19RCc<A9HRdY;43(5F
// Ee@3^NP6?KMBL0UeVCZa@A^STVU3>]75eX#c?fI^0<OQ\64(]Z\&>g:EFRFO67R&
// 9g=G5LRSQ-1J((9CBdc3F?ONU-3/7G,/V]]&ANUIVQcU-&L69;KZ6G&ULN)#WW(.
// [A7QWT-Z6#95-I//adcBS/W_.Ve_:91]IC_Z)EVe);Gc[0?PKKd9@>-GQ^fBV&NE
// ^6MHRX2:73\3=c9?f_RIfS<<_FWf,g0_+(bf,3dQB,]]BUB\^f>-UWK^bGWN^I4R
// Y(CPT(D#1f(7EW??C:83PAV(D4PSVa)\=-EJ/FGS84S[5MW(/4YDJ86H&+Lc=2G@
// DGKYS6CQ5QC?4(;BSV^+Y67I.V5SDCL8F,5UWLHI<YA49&<gHA[4TK8#><4II)?6
// 6[<-F;E63W2#+5>]C\I&Rf(:GX2WN9dZbDg8QT3NG@T[bJ&H0,38=L1ELS_2/65c
// M5(Nb8>I1aEG4;GJ)_11N3,KO+)EbW_(R<1;=_;15>1VKU]B?aFY7g-\K#0VZ&&g
// -gXeOZYdd5?)2[g.C3K&S5X>\dF0<<.)SN-ODa4T:_DZ84aZ)YEe[4JJF/1H4OBT
// U)F,0B(30BMX(b/F=V]Y+83UGcLMDfM-ZJ&8S+IAD2&([+;/ZSgFV+(b)Bb-C3H)
// fIa,SG.T&P^d<>JM?+8Tb[U9Y,AX/2H>@V#X@c+XN5I7Hb:C^]&8>B-148#(TWFd
// bW\=I/dFQ.&4@=cN-F&-<cKM7ESYKfdF>YC79<De(R1>(8(&B(G/K]9e[0[_.YB.
// M:f@=>bCE]2]W_M]0a+L_38B[2b-O-LOaEZbC9J28d+M^>?#T&DgdS?5a05#K&=F
// 13ITFf/GT.3[8[bXSO?Vg2bMCIP6023P-ZETT,3OLR5U31Td-Q&3X9\cKP&aW&<3
// VCL[S-/74GQgG[+K-@_-:K,B]0ROW(-LU#7Q#)DePb\8S40cMIdf@;&Bg4(?WPNg
// a-I71?[?&ZJ@I+KQ@FA[53IZO.0+AJC7Bb.A:+?=:FA2)XY2MOg+A#RM0;;gPTbS
// E((fbLF?Y,FN1a[#9G6CTNe(gG9CQ8OFBJE.R?P\K_/)D:MV&L)K?\W_8BYIPVZ2
// YJfXWH<YdD,T_]=5f^1,eBCf\&cf(2<2Q2FNDHC]X2)\KW_M)&Z^>ER([4CbC-0\
// @U/0_[(#]M@=N)><\NI+=]+=70Z:_ecG^K+RNGU;8+D^4e-8+A;<2e@UeNKe?M&Y
// VDK&X>PYTOBa46,&+EO5=@ge/e#GD#OUfaOK\<X820?YP&T:Ye)HN\P#R4Q+C0UT
// c]<E4QdCD7Z_6QONG/[]]_#-_TY53IE4Wf@.e22\2HDXQUMC13Qfc@;5M]+FW:4H
// >.)?]db.3).W9WRDU8+JJ(I4N)D5])&I/V_f9S#-bW.=\=gG]NWO:-49V0-[_KQ1
// 5NRY4(I#Qc^0@)e/-LDH,fKdR]7I>(KR8;Le58(4b\P+CN?<e0E=.[O9Q(Ya1YZN
// c@_ce<]R\7BQ#9CNO?TEGPZ_L@V4GZ[1TT0(LZ-R86IUANBT:G(8YYGBA((VBL6O
// Of2?-g6V.0HB?S_0<P+Q148ZRPN^Y?30;X1XGXA>?QRc9ESaUdKM[H4\=URMJ?cL
// ^D+#R+?]^e?B#Q>2U^a[A9U)06F70Y/->8IJB2VXVf@SaJSV[g9g>KB=L]O2:edg
// .+YNI;]WXI:/.a:G3L+YRe-Tdca@C5DM73#3Y\#Agd?T8WN(a-B]Ea\F)NB^IMMK
// bVcS7F/-QOOL&>=G=6E=(K.B8^4NH:HN@+CM=.8)L-5HO>-EDOfcO,Ba+aPW)[85
// a.G#64ZYA6N@AXgW^OSee2Z3Yf0b\<g[6XHMFHd0NONIGF8Ub#.1-B=>DP7?g7<a
// [&cJg)3FZO/)Y4IV.A.#YE_VL,VOGQIB#5g0D1^@<ITTf?aT/\2Q<>fO<VdgZJ:a
// -Q;-[M(eXC1C6LgD5&23?J./KbJa1\P4_g/gV-W4>DE?QB)_0TPaNYT\DID;.7ZF
// g\1ca_F]DHT,:)CYc^EG_)>-2a:N\4.HSaP-6HU7D&65XE3AYIUFc\US]ZgRYbR?
// B)P.f:.(K2U?Q,NLSG1HGJ,>/[;#S5RX#Ag]MgH#C=fcU78K?a)4V;T;eX\7f8()
// CGF&R.54OeeM9b\\;#.cHeUIKWNgd,+Oa^KBP(Y5]E\97:P[.f>.+-,@eE3?Q6J.
// (E6(W@WD/Z5G>G.G8e@KA8X/\^,#4B92[gg\d&S#&)Q;VF&(\?9_:ACeAa]X>,_^
// 5/,&F<HYeA5bHFI,L]>IU0E5LRCKbYcb)DFVF.+IOFgHX)(>._9V5.4U&[\LTa3(
// \6dd]C,LT6^)S[A[,&5TH2N9L5:C)W->)LZ+<&_9dJe(f>,L[J:>^Q63X(V>FYNX
// 42L>)LX.UF>M6[Z4?c2Z/E<a0GH3P<5Wa6V-aObA5/5#T&ZQ>)4YA^_>K0;D.D,C
// 5[7-X)bQ935g/M^Id_TW@-d.DXLQPI.90Gc@+?U0GY-HLDK;SW&Y[3Zc4W,Vg=#,
// .:,[,9-N/A5KA^RB[bBCAOM-(Fd1;Pa(B@F]>[__#-N9;OAK:FM@XT\Z,U3dZE7J
// f,KbEF6S)cdU<_3?a:0-7VUg:)BW#7RT7[5TE<I<//dS6b#W[Y(CI25IN<9E#8#c
// [f2Z#V^W?^X;.0>D4T7-6)bB^>f?_EN>]79P=<OT8^fBK,\A12^++,ANU--(,L>_
// WX/(NRH:FUB\aD7bH<aF6+H318+M^<.GH.5P8YVGRf3ROQGJ1e-J&]_CNX_01IBR
// dM3gKY^_R\ED,)-T\f^8<I@Ib)KWV:>C(MZVg>E<>EIRUDXee1IGOKE;3]+9ZS4d
// 47&JE[,DI(R29:0cAWMc#[.Ub>93.^5gU28+e/^KV^W(+@:>XVY+eJ_Z,&<L=514
// ae.#C9?@SgL7;AbS=/47Q)_dgF^KKea?8[X(FH<PB_F;AD5B;\(:RX#L6V,U+<:/
// a]^5[ScJ6-U)),E>3MC\d=1UO1#+(37d17;H5c39-9;W3]C^VX/SD=<eJaCMUJE>
// 2.-LfYT3>U[MRgbBP&GEEd6:5[,cEE.8H)H?DB/X+0I29ALH5J5ESdM<OZPF&7-N
// /N1KJ5MGHU.]C-760GBOW(R5[>\E:Y,UOQUfZ7Z&(e#PO_.ZNX3>FAP+>_&EMO:[
// [H3]D;R0[884\]bF1gb]DE2K2Q\>WC7>]/4LEYeX/@.KSO:XR8+#H]Oc#T,@eZK>
// ,7@ALSIf@d6@Y^^G1:XU0X=&>6U/I;ae@T7a(F6[fZ?2D>.=M+N(f8HE^T()W5Yd
// 6W26RQ9JM^#YXSCNQB[=4QY)N_?2MCA1cV@^8K)3PSDOOEe-?b-Bg\97N[O=:>fd
// H+UAPg>[KHC@&].3OaQJ3T^_0FT2,a0_\d3cNY@NF4KD9,5>6.+J\OJX7-FE;cd1
// .V?6/:-0HXVGB/,-3=,V3BfYG7[N/400+A?35gF#+P>gQLH-ES(\5BT[5OP6=WJ+
// ^N1#2MTV.a/K^._BPC<=3Y^Q1Hbe)6gdbUK]JKIJ<N&N@T[8U>.29#RQ6(Ic\OQ;
// I^2OHcR2K[?NP7B;f(\A=\I;3g8C^UQe[U>R.<b;&g624Oa_71@+ac+3G=+Ka=3E
// )N3@S40GJRIQ6:CSHK>=U07Q5fE+4](N>3e.cS82_N#[SV&HTF-W2AM<U5?NO0EZ
// C-6YI7(VJKXFKH8FEE]H=L;GN.G.I69;9OC,_Ig9>7A\\ZaO2;DEH_1(.HGG+a8K
// AJW/+R<NRBLAM@_OH)&@WW6)-#N_3Q6a2OE1/+DIa3NF\>T2_)B/Wa\85\LU+I,Z
// ;3+UJYLcE96HJZYZPEC5-P[BJ<IT(6,X.E>,GRA<L),@Ca[W]D\3I^T<8KYJ2AeV
// fIY\BOYDDQb<L;)Y:P;0W?-fG5#+@A=5Nf19/1@QDBY2UY_:,9H[0)P4N;1..)5N
// >/=_FI[ROb:AKb@>KL8b&,VcOaO<ODd(--M\gS.78VT.H4\Cg@UDN1S@Zg\Y0@Q6
// VMS9>OWR#TTbS;S7d)B?I=8LGeV:W14WW,[VR9&;II+bIId23Y2PP>1bZQ7AU5]1
// )Td-0Dbg,PcFQJQ@O4F&2I2bWdX)Pe7,fe6LT;b_BYdFK>/\P@_dd(IE[OUQ6G?^
// dF>GY=BY^AV6/,XS=X;0KfU;_CWP_,;LTA3W;0aM-1\=4[J7eL82Z3Y0K[-ADOYP
// Y1X6SLLC0\/(a\4S_=1YZD-RC,:(D=@[&Z=+:)3\FHDSbAYYdJQ-d:Y5@UXWER&,
// eXPg+3;eFd+HfX)RAXP[Q.^d_F#T2F\O791V\K(PY0:9MT9eU7G;fI[VC=2FJO\\
// +C&4,>P>be]4&+L\LeGD1R@;4d9/JK/e:WV#RU1D/AEKY[2J-D&#gWSdTV8YR-[[
// a)=7L8JB+7E)JgOR.BM9WF5Vb-E)YF;UO=<Q2ZeagK<8=RdDfcL=7(#4]PHKI-D(
// K1@A_gX.4FQe3BR^EJ80[47dD,?Kb4[2/AC&H)&Y+UG1fV2.L\bFO,)3L1STXa8T
// b(0V+Fb\<Q1\QX<gR(dWgTgE.8^M^Z^B&Y0+DNA&GBH=<7-c1[X<G:C9C?POSg=M
// -W+X1^GRNT<:@>ac[4BB9/#UbSIK=W./F6]J2MHN.cW&;X?62;-OGZP\b3H_OPC[
// :=2f+]e^67aWS8Be@ABR0(2N.I[OcdH2P2KT-+bDe3ReMV3a#5V>)]MUJ)9_CI.D
// BV0U20]F/+X8W9QVD(aTcZEMR7N_0:OY1O3M.BNR(AK-R]HRYEAbKC]Ye:,1B5?I
// QLRELaKIRG&3C960:K0OaI5+2<HFABMC.2[JV=b-G^O,/KN^[^c]e^WCD\[7YI:L
// 33@F^<cYP7fV60XX>d9E9Md,3L6?Z,b\RVR_X=cX:Z6c>_+e1R6dY;BT0VPa@XPR
// g>];3PZ,Le@RM06C?3Y-\LUE4/&@V_HAN#Y?LeOe/GgU#Q,>.f)/N8)/cE0UNB)1
// 0G+c3/2dg74#:07@8)XPTO>G@c&:3Z9:U9J(-b8C7[7<OK[D5SX]EHM7?bL2/7JZ
// W.)c=@N(4DP[[K(5([8V:8H1WF(9_KFL6)LWSZf30T6c<]WC.A\X-P)8D4T.F\M/
// >2==OcWaKe=\,O=1X,+UDRE4V&4O9P?_42YY]NOVb93)..[FGRXRYF9&&::D/B+g
// X9ZY-P;,;V_U+V92YN^4f<1@H4BWLH&Yf?:9+eG2dNZeDZBFbE>JF7JMaTORXY9C
// A_BIdDOQ_N/9[b_N98MR2CS7Q>8&2c\9W8U3^]]]6X[T6H0L3(fBK+-KXS9/=,HI
// MD38O9_Nb:f/8Q3?VLUP,OL>(7aL@?91;W<OHD&>.Y8bDT_99COgT361IJ5>^(T&
// U(CC;=511Q];X\(_?-+<:#R?5,&4CaA<3cHN\OHH3UN2cT0JM<JZLS@RB1T8(.c.
// DDU#0JWgRF3PY,=CKA5,9DU0>N?7]?D-f^EJcLGgJ?^6NT#CZ#d<f[WK^5M<]S=)
// c&(YKDF&O+-5H(]HaDSBScTMC.++V61OV42DKR1M(b11F_T5&?OVD9;>0OVc<OGc
// F<3g)7WSUZ6]UK>C\\_&3J@0TcH4_AK;4O.5-a7CA[L1FK=R<V[6d+Q=P,_=5gM.
// WDR>P<?LRLX/V],bDP#O?(,3,J;Y7EYWXadP6AFVef;(S75I=C/b2=gT3]>./-&S
// \gWg?+;_AYX(L)b5MHRB7;6@53(Z-C#JY>\K,IJ6a\_4+PHV7TQI3VPf/3#@Y+<0
// 0TMN&acQN.SF9K4T1)aMaRY0#69I63^4@UE^:1?RJGR?>&fJSg2dMV7)^3;8@W<S
// Zc/>>EfL;0c?&8b\fGa?_4=BVMIbL.3a9a>14dG]L-7:J]14XDaOEEgfdP6N8F]<
// .D^W].0=KK>aNCgB&;Eb=f3=SJ>_8>DQ6WMS\AD=5TaCR7[#[cU7Z_AL.W@T@=\8
// _9?QL4F+=+XBJV(8.BGKLZa?<(g^6BECd8ROTF9W.\Z-B>F8=ABAE2PTdJ_[461a
// VU;,8(3#[a9QE+Z#_I8C;4(Z1JOPDJR&C0YdV&gV1M&dQ(1_-](YERX<O2g?JfX;
// #?LHMI^.8A4L8g(7I3C/P>H)_e.K1D.bT<LDS-#:70UfbZU/;6K#4BU7X9c[>JT9
// @)3ZO6U#CYf?3a#43.#S#)e[P<\9(X(Cd7e7,1ZY+F0.4Q,/abCOXE0#ccN70KT9
// W9/;=QDJK.10HcAC^7(AHQ]g,SEPNG:>b.UE1,_X/DG9^=PXN9#T)LB,PT82I7()
// H60WGQ.YDZG;FBHg6;G/[(NQP@FVZeLF>f=(Y3MLZC78P^/-:SP6(O]IN;cgc3V(
// 7.RQC=06g-(4))I3R\N(M0DS;].CN0@dU>=4I/2:G<_Ac/d)aBQV+M_3H:PUCPW0
// Q,Aa2QM7MDP74?dG7Hd(BG[LXUY4<B]^IXW9FCOV\WRR5PMg5ad?#IB2W79D#IfQ
// 9abO<c&^B,@BDFM2U\.a5)1IQ7(e#?#;</;3C+-X0-TR]XYC:+U@7-bDg#E=WUT-
// 51X:#NR]Y;c3f?cV;D\Y.GU-62VJ9.;931bbQ(+eHdRO=>LQPX6-;P6<0(EdZ(X9
// C1C4Y]QPJ795I0.7U=CDOB4g58T5TOM1.&Wa_:QBQAbWge6\=73X13a^=PHW^<5E
// Ff+KI_@Z[a];4dJ2PHA@9S3?LECWRe<#,2-9f75&&ZRC57;QDZIW.(FIV?:+:)CF
// =A>A.C@[dHH8gV@(G<P,)#?<;J)ffI@d6Je7;HG8X.A>(RH]NOW?,MdT<B1cDXf8
// 7^/LL2YF2H[A(L@XdB8;2aD#eHFYS<&,Wc4U&F3H2gD0,Z@B?@e1Z.KE)V1UI?gg
// 6?W0<g88FdcD5LWN_,@^]8((+<fL@_5N[\(^IP?;EMTBX;5MN;4-0<(NWSBg#aF=
// &:H;_W#ec,F9]e#V?a+7/)W-fKRO=E3+Z4HFbQJVR[agB;/69Z&7eMO/,If0\XI-
// :Hd9cTUZH[V6Zfb/Z.-<-L7;\#He,4)V:[bAJBHUeB#N50&N2L&CN(K=ESDJY_LD
// L/)Y7A2\U6G4290V5(_PCT3:_S4]aFHVN@a[?C65Oggb6HVC\c#U,MC_?BKf/,TK
// gJ^[5/=@d_J.4.>?;U>M(V>_L&F<&;gL0=eCIKW^VM2W[(dfTWe3U=fU/59D_,\I
// XC?V]:M+&.d+NBR^#@Gf<b8RY5&:N[G5ce2J872G1NED]V\C&&16W66DQfNgM,)f
// aF\(KK\7f@7C[9/f,PV;E4J/bZ^(O#]-Eg.?JB(1Rd=,fX<feYb5K^N;&5[QS6G:
// 0[a[-=)aU&L?_KJKIREcIAbJb7HM-17OUa.S,1fVEG?CGMWZJQQ^A>_?>gAR]<7T
// 3DA/?_,RA(c2)GaVMc:JMH+bbAa9PRDbGa[_d0J;/9A>[CHW8KfL0H\S3EH:XX]+
// ?.;:H7B:Q]U&b.Z)Z?(XKD\:MG:[dZZI+CJ^JO::#-->.+UF3:.E/F&AL4^,(.X6
// H)1O9F-\/Y?XHXg));;BSN328/J5XF>Q9R/?V2[1@4@)T&]AfLSg5&#^Xe(.,V-X
// Aa^Se/Q867?G<e0[K>6?:EdN;U+OA-H9I02?C.B/Y(EF)<O&+IY469Z.NE2[?DPX
// -8Tg/ZPgZ^ZNaMHLe1A#R9)9G/@4?AAUfX4K;JFEaUD9CIa:dEJedQ>BKK\1SXV1
// G^]HF]TWA:]&>(R4YNGeN<W+;5?(c&]1+E8A]-_C/UbPHcBNaCQ1REc-1M1,K.-,
// EYN69YO\c7&W3)<_A\9B;,HVTTY2O(;cL1+[)_eLUO@(]S>RB?YD9WgEg0e?>cVC
// 20RaE9BG65(_U??B@&CZ&QYJ,B)DJUDU>GCb2>Z+87c0)]0+Y4a753N0MaT,/AeM
// L#6^JRY5M0]&V2PCR],_:6^[I@;XfQ6I(-1K(?ZN7+MH15-R6TN-PG@eM\;.S6Ib
// 4J&XYO5M#,fe-?4I:ZF+HNUO@4bE;(/P.1,Sc-]6c9:7?8508273W#PJBMM9:FUL
// 1RGJSC,T_CMR&6EU9KYb<<:eUU>&5E:LFWX.<0dH/21K2(.Nc1Bf7,SE09b)@QR?
// V4##]bPb2IP8gRcP_U)_8&=Z7IM1@A]bOaaD)M8C/:<-0=M4Y&M/8E6-0]AZg>O2
// =CcQ<J2VI\e(/:Qd#<[Y]?40W1E\AH1a>g6[S_ZHf,T>[R&(b8\H;9RZfg@T.G]H
// B,W/:EWPUI^+9O2-D<2NPJa+FQ/:U)@#9N92MKD)a<_Q,<Q2YQ;5Y]EO:aRM@GdT
// UP:BG_S=.E-G>P4F.YP_XVT3CE66MPF/SU8cL>JRN[aW=+5>>86((F:]8#?U9,<Q
// /?D(SXQ_1Pbga]fK8X#M9]c5>.>YgLHROabU5MLVS#<2<+>HLV::O;)WFR/A;V5?
// fe0<U8[.4f)&[_YV9E6B(J>((K@C8B-/MD>8[P)&]>L&f:(/:A]FdXIfD]F3KOBL
// IZ4ScAF&6>S^[+SO)?Sc7eS4)+eH1fS@EX]^5P6N,3&022T[S???VH@R7.]/L+F.
// J6bN4P-=?CL#1Z:9W?fITIDMVXV;M7@JU:cS@RG2I?M0V.RG?],HTPbYa/db+fXE
// Y\b@7B9:bf=#0R&^<),:88bGI_,Z6&-:bMJY8Qe3KB<=W(I+_gON5I_[6<^Y)a)A
// FbTT438\)[=WAD-a^I8&)6?,P@5O1QHA32P6d28O.B4L_b3C;U18HUJZ(O:O+^OU
// .B?G[O(<W9Y0)T1OYVZ8:E_9fNR1>f3]9QO)+MWbKIYAK1Z0be+Y^FKSGI,AABUV
// 6G-X=B0D)AdSZf86f.a&LC_C8K:PMS^IDPUc#&A6D;eDGSdP3bR,FT4QW?SfP>\1
// ,C+&gOecG5R6,VVa\Vf^C_R(bX\H]?ML0W-2ZD9]g-[X[fVKRc(VU^YH9P7UQOLO
// FPL:RfEWWLBMVL4&G+6?I^_0FTf\CR(Ge.7Q6<58BE2dV+[?\eUM(6H?:V7+C]_V
// \PO?=aEP(3NFD1OZ9>JM)D&LGU#79d@_4:(4U^Z@T8cQGR(]\A<V18D?XWUd9CCB
// O7bZPS6P,ZOR2cK@Zd<@VOX-KXZU9<;4TW1bO[MX6C@,BI5D:0MSZ??9+c@+N?F\
// <+@Z+-]WPD(-.5/BR3Ceb1+_<B(N8Nd_5+J:d0RF(fGd8FV[&W=5?gPD;2A/eKBV
// Q[:I@C^O:\D.U<M^ZN68H[IS<44Va:\3&-[;#^_8328:OFBH/5c]eT.DCJE]]3>Q
// -L9Y#-1S:2<R?Ba=<b<=aM)QN8b5K8T1T,S0d(G5&f5(0T]N66TRA#g5^;X\>7cD
// YDgeYXO0ERT\E:G>;FY8=ZM<^_O2[&04A#BAae&I>]Q&BTAGgPI5HFS^e=?.d(>)
// R25B>AdKHeH4N4aMd).d3;M0bYSTX]-3[e&K<4=)@(47O;<30Z^V3U;9CB]M#1LI
// -(0C=gYSMC1FY3S4GS3YU_42ff(S(RK?&74\V7D^#X;XgK)M<VJV+06;NJ<U5=O8
// VIfXGcda/Ag.A/1G;LEd?Tf\G1BEQLKO?<57)7[7g:/F0RIRH5RX]g4^LIV4WMbR
// @R83F_]-Cg#]NZ:a<JA<[d8Sf3#(-8H;R/?#4BD)&D(FGOS3aS=T@AYI7OX@RTZ\
// ITbS[Qd8AMD@)XD)Z+5MeV3NCa:]ZV7CU-)M>WR95I@+,8AHeJb;U+60#f#e-\4J
// A.UU#0dQe9&0dM&@+J,HN6Q=^A?X#CdP9T1D604S0::SeR<&;94eQ?TZ=1?G5_TI
// [[_;?D;eRgK9^<Q2F<OGL1=.cY8&LX[(A_/d+L?0RPP,7P)S6/H7W@\;0HBb]VaK
// :2W/]?>+=XCC-&R&8T/gNJc]=eVN88R1XX#gT7C()FBI5_b]JVD@Je\>,3ATE0]2
// XG2X3;EZ1@6S;]J=e,7LCVb7Jae9]W3@LNeBIY7,?gWO4eJ]><+cNB/BLS(]^FXb
// Ca>=5-M)\XEK-b&GR^O45IHVE&OP>&2KNdJY^#DNXY;HB9Yf+f3S6XIaAGg-56AQ
// f1c85,7U;90D=aF.HAIVfJWH4.EIC+YG5(7@=NaXQe]#MB[.QUZ2N:[@9M5)/6CU
// K13/8(+P/c<bLF>C<#b=PR^a^C=8;?3<^eR5[db.6Z&,C>)&46OR6F+#V1<g]JQ-
// [Q@.4,JSET^A+?=A7N+\>RT&/5:B0>F:bGf#BL:eaW+5LK@BOAO>/Q<,MKN+IT68
// @d@))REIZQg7&CWI^6N_L4/cGfX8TSTd@N>GZb<>JVTA]f]f@_Z9Z;O4<WF#7DG^
// )cbVMM\74[]f:E:4+cfF@>+V6+_Q1CSL>_gcZ;J#0Lc],]#AVLaG2HV?<LG#7IfF
// M\0cQ=bRW--P8.D2K;TD(9I7d?IS]:gUB,\OZTD(B2bb:JN(NIK[/1&2-9,db.Of
// S([U#TB5aI+I@d=KN)>R.7cO(P8[I80F6Kf-<[(-Eg4\MHb^.?#VB,[?S&]G6,C=
// +O/H:MVTMcKL[-_VgW\&Y.g#bBAcY68Aa]Q:VIQCSc<e0DP(c+7F>V6Ba[OdQfC\
// >XX\W-D=BWcL-_->-70)L1,1.63U9DbH::4M.?KOG,8U:@W(8B02a;Ie8Md2?BY0
// <,J9\R:6?35F:IZf0aZ2^efYPfda=P;Q=d.CgeJXC<XIV]CT.LFgI<3C=3PF3K,-
// @B#SQ3f[0fW&I6]:e>51UT&e5&&Bd?Jf84CB=aF:&9]cJ==)OS(,QPgC5W8cb@Y@
// G,.b12g&#OFBY&QXgB@ae>:-=V-//[&<75[fPFLXA8b032f^gW0c4A9N)@UAaGB[
// NIGVa2S5TJ7@_c0<?fKFID6(;0b2(cCaB&Q<T2A9Q1.P51d@C.,e+@/.NBH9B-DU
// <f<#CJgaW>&IHD#G?Db8U/R&Q<=5Mfd13dF1.BD);<E\]G=\[YMOF3gbZ:/)\XO?
// 3^AJ)225J?BXFZP0e=)&VW&#SCMIC>O3[F=/EBS99^SZELDCQ@=ZVF:>U7@51OC<
// LR.U)RKUC/)G)H\?#[^_>G3DQFBL^bTH8GEH4Y0#.X0&XTI8GXGYD3NEfRIRWR\+
// (F]f[#I<:NM/[ePQ2P8B0;BH@]IgA+IPK+-QMZ<;Ue.Lb\KE4XS:aMe2Y[@McMP0
// Ff+HD/ZWb;I&O+(XD:;<_S8L,P2B;#_ZS7E<Q6bG_?EU85Ee4)<[_2X_J&R1g:/;
// c(0M&QIg7]28dBe]TIQ3AM8L#6A1ce^?Q2>W1S@U2)3d.C>J9J&BJQNZAdA([fFI
// ..UFb,7?)-KQ]g36fS,fKb;]Fc=_Z4Jg@QL3MRB23Y>PeXTaXCVQ&@Bg9X/YYBFa
// H>9G>[/:C56.+94F#GeO=)X7S8T67SGLIRJIX_>]8=&#8eL44V3C+f8Q)&-R^#=V
// cKZ;>7:8.IGg<DUc(DYQd61_/)+YP>I.+A\C,0>5@#(/;1&[T@9fb0,I-><TfP-S
// UJNB2_PeL]VOGL-D?NQ1);X>TU^U_W<:T_@[ZU12@#1UKTTAZ<U<W6A1Q/KM4d[9
// a5bV1c?=^P9L2A;H5B16a@gVc54H33AKbPD@N#:3A.Td?7KCL\XW_8<IDc#g@0N6
// I3E]P^40:43<>.e8:5,LI>)dX)#-We7fIYQH),X;DH23-QEK<;/<ObZ.]9VNIcBF
// @RaX3Z,EV,W=?#&/TOA]]IX\4SVI(YeVTHSPO5+J>PL615AW[/JOI=BOE#03#@+J
// N<OOdJ8Ma]>@DPAWd6:J==W:W2OR5XZ8<XI^EN6U#e/EYSP3225TF[2dQObSef-]
// PELA5]95b3dHKH=LP?&P9]bOR&TE9TMV_/a=a+^TY8Z+=(86_25cMFHGW@+J),Jg
// Pb[&fcH?TZ8Rad67b->Y2TdfA^c1,C/:g=BJZ>6cIC^E7.N/74EOE:D6FB1C;)O[
// <,1R7_<>B>)HZYg_3\bEEKd,<UA6DSE8J<.NN^5EJ&O)&A\OJgKL^;^a/\8Y>>H:
// &02V4/#F<8FL;M,V+=^Q:>,,W]ET5a@UD[?HJ>LfSD.XUAVd]C/@NY>_R7]Pf.?4
// (V]<LAgX]#Z+Z45P(ST6S7)aHa.c<A7b#-1K=\WZac2Y/<UZM?L6TX2HIa[>:N1+
// (#^7.-Ob>g@MB#WJ-IPCPBA)J8]R6AJ-O8.e.[/C<15a/3;D3XWOW,BeSPQ[O-TH
// KI@R2O1?3-?dA740]\P.3[_gSECeA2#7g3TZ7F-6152Q#c4]0>HWTCfKdM\66H72
// LR8G0;@R;@>_5>)#:JRc_]V]7<5g#LQ9(BTK_T=c8+d5R-42O3K(fK,SfZV_O:A\
// U/&/CTS4JPYc;GA(^8/GMXVA\=,>BAU,UH7JT[#bSLQ,6)@VG4_W&-=:_@4f)#)H
// P.gJZ4FPWUd-a7X:)\g<T1.H5Q4O,&PL2CeWZd9-V2[:E>DNed)e\_ZHW[HIO0_c
// SMS:/@,^5:UeU^7;W]4e,gF[McFYG]ZU_OOB7RCWF:AB(9LH/C=8W.E(I49?KTE&
// NZ<AVcb=-\O?,gF)XEa/B8(g#+NR,d9b+ZdAU>\@I4\c4<_EN_8^5Q),RO4,-P&H
// ^^?]aPCMf8+2Qa\]e_=#.C74b7Y\>-eE)R@N;U5?<[1-G\JH]HPH(3T6(OE9A4fH
// 3eI>B,Pf0WEc4HOIcD;D[IaVc;Y5d-K(RQ#K^H0^DN8,:?L>?T.H\CC[-3+R175?
// D3c8B:dAP8-NB]3a(>S;6WQ#HY2f(67CcfBde:XZGf2eaD]458D+-(G.)8W[A1Zb
// #;1VIN+d_A^3[ER01bg\<b]T:,>F78dY@_SIO-,Sff/75b,fI8:O5\dY1:B)O\J=
// 2C<Oa.8d]AXPbFe</98=9O:SS@-1Mf4PbWCEB3D3Qa5@S[.6XH6:0a<1J,XAN<@1
// _1CMAXSZ<DHV9Na/L;RVc<1UZ8OS6^@TNR:NA[?+@fbgNA\/aC>XG<WKD@1^E59X
// dX:/YDIT(f(]E_;@W=SDRaNS@9_-aVIJQbFXKd(;&/bH>#dfDR21\fA&>430&.HG
// 2I-_=.^Z3JJ;=d,PYCcCb[(NY:4\[[#N,V(0,0_\H6,(4YXV[6H<II(^)D7G8f0#
// AV:_5/a;/g)\<P4c:MMJ>gVcL&2b>Z.&I5<#TETXVc,@J&@.\4cGVWZf[3A6/+[6
// 2Z=]APZf+:9ZcGTZfSKVgS^<EKC47a#RW08/9).[ALbV/-d6MgB,32a(d.?HPCM#
// ;4ZDEUa&<D>ZbeVg;Z44c[&.7N8RCW<UKB36N&>),Ff_C#0\Nab?Jf::N?fZ>e;K
// ROY-.)H19RA+2g2BBGG)&/+BC9@\SGT9T[LO2R/\;U3?3._2;TP;3PXcLJ,&6+A@
// (V;_-c5=7ND6?=b9+3/_IG)T@^0GI-H89+J-G\4HfZ.e[A_d/+RbgC]&F#U:V2,a
// 0IN-)E/=cIbGSWfcS9Y@-A,R?:e<A^02CU\Xf0H13PJRR#T9GI;7[;2)+a)<B5/2
// GLb_gSX7:UDZ#b,W#W/0ee,X_--TDH^S&A6<5&J_,/&ACPgg[3_M@ZU0CZ_G+L[N
// ,B<bM@#VVd<\Vg-SZ?eKX6Zd/NNNg=#G)fE#g:7X#@@5LY7XH=ZCg8)POXd=,JX)
// P=->G_g:GHG>[,?cR)>VfD>\DgHVC<6.HX=/eYgGIb=#fG<UVfSYGRcC0X?1[;S7
// HY#TSMNQe5R+a04/QgDKW2SMQ703V(Kae/E^R7NK)3W/4&a:fES)?C1AZ3-9AO=@
// <6S0:2RFTCXa=&,:H52,?_f/^EBC]5LPe<CF3aJe90+8=7@d)>[\RATeEL:J^MOC
// ZQ=XcG]b]\.eb>0:ZOQ<5fWSYLc2J5gQ_U(\YEaJL]W<AVB8&:<;7e5YG-#967/d
// 8F.-&7E6D8HL/KXV=gaZf^eQ;6OX+QL.X[#B^FDZ)M8J?/J5@1Z<a,IE-RTE_O](
// I.LH0LYW]6BI_8Q<;.47PVZJWG17V3TeE#ZOMJNK<56O&)c-)4=R8S/Xf(58PR.6
// G\bPf5R0^]1F5:ZBE+0e\K\DQRFT.97@:61H00+U_#a1(CA:7Lf&g5:8NB7dJ8.V
// g8S2SJD((@)cD6W.V:bA;[__3Zf:VLSH=BH86e<+3g=:aYbT>)2HZLXJ/RQ29G,[
// 43.Q0&/FRf[e8ZaNB3</]<[]@&d87ZH/37S6@[1FGCXd_]<CZ=X:E);[GfES+Y@e
// g#gb)>K1gaBH_L1FA/Mc>O1J0#3\UK54M+V_&I3N8(K,JZL=HB@8>V>CAJcN?9SP
// L3P,B[A?-GLQ8V^+RHc(bZ_1^gg;4T.g]_RBZPTD:03fYaPUXZ.@4(Re?DbKL)\<
// acF>M3&+]/3AD6f4@.b=YJ(/7KF)ccT24;?BF3\G_/:g:#J^U(Hf/T5M&)E&W5W.
// 3QN>(7>Q:L^Fd^NDF49T2C3;aa+XUQabXD?45\XRa9F[WQ+0\=aYBDR0,0D,2^#f
// Sc>S/1/B\L^P/)41Cc2@]<Mb9H[6d#&ZACa_C#eB,DXZSX1/_fgDG)XBZFg?K&9D
// (\.GY,H7\F(CVBcU?14g29/-6HVOLce;4+?)&SEVSQG3/YgE)?6aC+?_OIU0Y^L+
// ;U@\C]@[A),DOV>A7QL53Q6]153a0G<]32KXOP;+AW9a??5BVQCQ=Gf^\c\UW6\R
// K-)267Q=E>Ybc>_+IQM4)aH<(V.]U8#9K[Z[,LH=Pe>X(=d;SEXDMTVU]Q)Y6A92
// cH)H+IRf0JgW,BA\:XaXCQWDIW]Zb7IQ)(YQ17KJ1e(caV3>&LW0B>Q&^U:G.BTE
// OYN=YG6DZ#UAGZ9^T]Z?:]?,WU#_^9#QeYY?LdEe\de[?fa.#dYBG_/Y0^@Vd;),
// ;-U>C.Lg)MV6U-@>KQVT.eXL:BW8+g?5_ePG8.f\K(a(1/ASO/FD1:\FU6J)c]IP
// ffYSgDAQ_]9&^BdOK_-RIG8S>.I.:8dc)R:]eH3ZGT2(edS,?;)\5a:6S:b-ccgA
// d#A=f3VQ.T&0<42aFYB4K>HEIQ7@[VY#G+VYH1W3S[MKGFG4C\<ddWS#VbB&F+a^
// ;gbKJSf;C]#/6\B5bRZTJ]7,A(d-Kd4:DabT1P9\U7YE]GEdfEaT@&MF=2_@eN\U
// SGcYf^7g)O;e:+g\c&GXX_^8gMS8VcGGE3[FfLS2Ng-J]QWH#NR^c.N-ICN2TSQ7
// +H,;Z#F,=aI++AUU_64cZIN(<=[CF4<X6IL69,J[>7R,JI+3DA&,fNXTg_e4YGX6
// dG:[15-AR-D:,&&STfJVZJIKKE+.3,SHY0T<J?#bB7YJ3-c)eS\F6aGPTR0\.]=g
// WAK7PQ-4^2,<ULO3ZOB8MVZJ)0(R7N56[BR+B<X)e)2?Xf\P1)\[,)0L62TM^>-<
// IU:IW)Y)=H3V9[54BU,N;/KP\^@E.7F)b4]]95H8Qgf)&5Y06K,XHMYZ)fRV,SKJ
// 5cf=:dNJ=Q8\K8V:7JQ[4T^,]ZA08dgO,R@ecT#V0MRgVA;OEU\eU7/GFS;WV56=
// 44.7Q7X:3[dWUV>[I\=SGG0@Z:REJ0^c)UAf;<a7[S+&\)4,P(#MP&1N9.F[82/8
// HV)]f01#d\R<HB_.6>N,[_0F6W@KJ2=_H-_,\YK;\G62OK/[GUUGc23W.AU7HbM]
// (@Ke+I>@)_?\5=GP[^[?F:-W+K((HT[;Q6bKZ/)6,4E@7V4Xf_RSa92C^GQ:Y>,H
// YO1ZF;PIeXf2b8,(VN>>1)1^6T#X9&e7@R-1HE&8M?cC+L[fH89R&S<1Q[IEEHN+
// 01E5d2F\WHY&]Fe2XO5-K2AOH0D(#B280g3R0WM@]>R<&^U15Z(XJ/H?HPCee,G&
// (WS52c6>M0dV:WeS;W5#/OP1M&]#9=\]34@Z7Q;,0dSLPc:e[:/c9=>QR1H/f1/@
// MU2NWTYM+&L/EL]dJcW^146AS0[#aF2@(cdSR8AB+YfCL=4F,[5OOab.BE099F5g
// #HG_]gCg_)\eK2YQE7>L9OL^Y>O3>0Me<(8R1K:>VTZ9_+.\A;8<&aSGH&OdLLT5
// (a9Wd[.7c^b&dLH#P\3)b8VSS@MXd^WE>PLQ<1fBf].)14([fLEdA(EF9D[DZ<N[
// 0/DR,G):/gCV4ggCQ>eC-YL>-cbAO-TYeQY-/Q.eZ#I7A<_ZNTOZAR@a\d7eT&E\
// Jg_E2#-<?dT<B07HfS=#Of.@X3B.0ASaZ:BdS=-)8;0S.^X1FDLLZV4QZ[=Ug(&c
// L2U?9YJ5e+S,=H.VZd_]00EO;F7Ug92Z/PI@D1^5]A;c0[Y-&.6BLT1GHLT7CI0b
// ]WHA<SD9Y5YV[5GO-fg_B.)7]:3=#SK@AM@Fe(R?7_a\(XA@7]Y1\fBRZY/SG,Q4
// \E](X\2:L@?4/?R88)6,IbcQDEc<eKY</._AeVf[&O]7bZ[aY1^,1J,dA6@9CL]A
// ^JYeXB-Y\PU>^-:7@WZU]XAI==F;eV:G,YC1TY?L2BVLb2-YLS\+LH@DCX_]-bdS
// 0/+g\+-#MRK)]J^(&[M-GO7]XcUKBZ2^@,G7;G;eIf/P)YR5c:HH([JE#T?B-,KQ
// F4__A>N:<&+JD#(YQCa0.Z[_g)@M1333cdE])]0^?6Y[.84f\]^-9=/N+?MZ-5G@
// .8)C73._98[:/?S5&??[Y-B&#V9O/MEM;8ZV.K_AVNc4DCZag2X:_2,R83.Ce/eb
// SBMf]43H(X<^Hf3#Rg1L\SIQ)>QHbVS2#1PNO?a1McK^aZ+#15;J,_b/AQ/@\<[6
// 8F++TN:)PGYPLJXFU:a4-c:OYBUB[Q/8>Fa8K>G&_4g?V9IBR&&/?-SI(>63J<)M
// >]aJ\M=M?+=/FMXWC_Y&f+E+4]NU,=&2H,;eXEbcM4_[&/+3e)#K;RU8^0YfS5W6
// 5X1fc1V3dY,M,\1-eGIC@XO@.JNN]#=EC(\W8J>.(&-gQdI6]&X.ZWb2XaS<X6FT
// G\>09/)BT[[AP1\6)1^H?Ud^T?<=UI6&QXQ,QG\\&0dLA1T/?R5,KC_2V[bP(9aI
// CH)&(WCN68L0,eMA(eF3FP)P#e4@]=36?R2/K^3Ca+BZgE=#Db=9a>-[-4V^/O]N
// #G:XZ^NS\Vc\S6U_SeLPa7b2VIJ1TW,1WXV6GS&+e-I>ZbN>4CV;&CS].579\6aP
// ?I83^g/DEPOE&<YX3RW7bEHSfDW)2<+)I[c-,+[d_#)eW\.TMI&[[L+^@P@+5[:M
// GX>TH=Sce[@&f(bWI_;=7KDKL5V(5H)a2@/UcVG\HE&AECJ5&-5=&8J6>LV&,Zc0
// aE@I[&6@HYdNdf8]CfCA)\NAHcaE7LSe5#FZT<DTaC.fFg1&KQXZAZGOJT]#@;I1
// 5b<(E,DDB4VAF\G@AC,;/Ne<JA@9Ga34,_cC/C.VN?g.Z:0I\55eR1_1]X?OP\d-
// b0b<:IO:TQNf;fPV4G(SDZ=6/gAUB&>Q[-\8eRZAKaR,YZ+Ag4?gQ\/7MY[\FO0X
// J2ZT/C1^E8JS/f6-5c5C5,&d0[LVIW,9@7O3QY1W@Zg=8^.ed8+59K)SB,K44.DY
// IUWN(O=#?G(14B]@=T&2/?N/Q0Z<a,ALP5)9Y;LW75&X,O=\?X]X4?/7Ya4(D\MY
// =A<UHA;DU^^HaU169Gc[-/6M#/]BQ2UXG3g9]bd+I\LBbG+D]Dg[<>R=<6M+OMLC
// HV]<ZB&EC9.\]c]31HTb7O<R5e^>ePMcK&Y72OEYV8HM=P(#6Qd2I3<edB,0RO.-
// J>Ia&&656C+<NDP[0_.8RJJ_YLO_)MB#5a:&\-MKFcYe08.G12)>E;_/X=A0b&3_
// <P.cIDg3.T4T1e<3g^1+VeB6ddTS[VATg]d#?#,b16ST0e=CG34LVN;E/);QRQ&N
// FFgHaXB(=&Q.@,\^#)^FBYc(f6&C?OL/RNc0@g/)-[DN;UETNWT7MA<RdT6\;@-G
// =JRJ3M5-4gPGBR)[ZGLF-,&VgI^4e->8-KK<)B>&Y1G.8O>)&0VV4RbQPC7Z2LG8
// #97]2_fSIXZYBcBP5/D\HGbYFEC\J8>GHZ2]ZBDC&PQ0Ke-.T(9Oc^(,PA5b2N>T
// ^Y)A6(LC?1;;+H0M6K8#5dLLe:WY6dAW[IG#?9DRMQGGK>7<Rd)PS/:Q.242DVK=
// 3FETF8/ef5Wb-gK=&e=3ObL8:,51/>Ve1AP79PcWe67)I;+0UTHIQe18/ON[,E&Y
// &+(8T+dcSC6I6ZU:PA>&a_80]ZQIe73ZN3ZGW2FRfF--E5E_<&<g2aKZIZ-8@-d6
// AG=:BOY8b,];S??g=FMYN?8;,EgSNYTP(ZEfBGdQf-6_S:L2\K6JCb4(2FaSG^WL
// _(Yd[SJLMD=G-ME-+QX<?XQWJ\Z^gR^4NN6E[YGJI9-U^1[5QPX)_ISg)F;N5@)/
// K9f(6HPf0S]@_]&MKcE88((#9\WGQ#;XDVO6[@fd>7WgUMP]NKRH8@-MIV]?58TV
// Z30g-QSeXGZBPJA1Qa>Z@41=2T&/;8S8SSUODBS_eNVI<MY0#N72>GAD/=K:XM/I
// aGS235N4_/WW?YRC6-:[<5.aRL\3E/J?ab\5.CI#0_3cHZ@.g;Z6Q9GW1&4?Bdd0
// cDOb3aF21FOY^:SI-KZ@S@B_7(J^VY#>=c)YDf=->N^e,5gQOY2WL;WQCae_PcaQ
// )g0>RgU31=b@W3^+&Z3,UAN4R85OJ,.MF0eWF[W:.JR@FDBMZJE^3YOUQHVY(_X1
// g>E;>R#I[PAbIQ61+B6^5S)E?aJ2RP/8D[,1S(<N&g<DM1N5K?9:@)33^)[e-W,^
// .W&6>cY09B,ORUOLdJ@HSP0bLVW6&EDJC+/ZeY>ca<\91\I&4VcRA/R2(3W68gSK
// @:+D42K[F.>bD:3bW(Q/.c0UgNQ75I=:]H_&^B;-((K-N.^D6c;-=P9bcT#NQKVS
// ?HX,SS9@+1Y3:XOR#0(BdPf+cS@&4GZb=>NB8M<7DRI(^KG[GL5/UE)\^/UL/0[4
// 507e).@.[5-?AgCOJ0GI63^e2VQY?gQgMRYNF7)3a&FAQ_7d?H-Y0SUZ)J1TAL(G
// AH\XaX6?aAYV3:?IS#dZdg#TU0,.8+-Zf?3N7P1g<#+D0;Zg14.1M=8^#[HAgR3_
// <HDM3T&:MeTeTdU=UI(77;8A#,e88._Q1[:I^/^^d]9[HLXaR#@0.W-f5^3\F,cB
// HZAO@#9CSab5\Zd<+I#HE7DELQ;>(YST_8^_35Vef4V+,:IG@BU?dZU-SSc\#1-:
// =FV/&fXa@B^4[6YD[-e7GDWJ8BZZALf?d=L<G)5cM>?Y.L@WORJ64[/:ad1Wb0X5
// 8>bIKZAN<FC>.X/<ZR21ELe:B)g;eb#4J/CVYe?#/U9E3,9P_N7D^DZ6>a:gN5Nb
// @<f^^F?(W3N[PfCR(.;;Q/;YM\UD[8#A0E^6Y7,d59#&.2=TgUb6/ZEOC96)8XE/
// S3OJM6A&4SSCgS3=HG+-.YNUNKaZV3_++dKPUQQZB,&d5B)NIQDR:<[Z7]:,XC@c
// BaW]A];_KH[dSc,;+FJ)>;[UBQ]3<K+0?8=Q8ZF(aAS=]E9BG96O2WG>TR8T&9#J
// YHDCD.;&R(9\D]c>>U/6L,UHDY@4f]7O)V3.6?6WMM-7=43H<V0WDW1.9L)5f-/?
// d=X/;CC9@L4P,YYQ>c&4McSG=S;@2XEL0;Q#bH.;B@dOCRPG?T;a<Cd1JC3geVgP
// Y(@A==&GV@8a#V<157LW/a^?7RL)=g+AbVY6d+:]0#I<#EUe&4)eLPL/f50PZS=>
// (YI[+JLg33U>XUREWdM5U2,@,+HE]NR#Yc;[C=OCL+WdgF1c)6AQ(g5J3F2?P-V;
// O(ZO#P]RJ.d^17.U+P1XY>-e127^SYEYP0_;)/&F63[T?_T88_S_OI?dLY)5NB/A
// YCU6IVIVDSSY39Xg,[AI8]&H1C4^+].00UOOGK#bg>FI#0D1KY;IYIOVO9(<@J0C
// R:cSgC8/.S,N^2IGC]KMCb65BcZIScXGePU4;JD@Me/+[-I^>J<.IH^ZVK8.a(\K
// 5[K&TYe/HX^OEcN]R+_2S_1EJe5(6\+>?eCN-R[I5QFF-S,8a06b7XdQC;C-/5=9
// /SOZP>M2>3d@OY+Z0_Qe@Z_?a1WTUZJ;55F124=<;I_1fSMdK=&,\cAY#XX9RPF;
// )@,8DPe_Q[_-c<MV&J>TO9&&-b>M18&UO7L=\A)\)c&;XI4>:8#5:5Zda7B#A.^J
// LXKSS78G#b6J]g@\VM?#54&;C.L<9?X6LAUOMbEX<FD_]0[&</53(@/;)HW+DDMQ
// R<bc\LYAL0NeRH.NcV#JeVGNHgHG3Z-T9e0]a->0Ecf#2V<)GE]MZb9.EP6O]0TM
// gfO;1=796O]a9AMY_5Y/BA=Q9G(Mf.NQ)>\T74E&e:O>EC8.,;[7W_.N7=JQd=YC
// ]QR?73<W@AR#U:bZbZBWA8@EH76b8]E@]7OKRdS>X>FP56IHDMa--QULaK_Ygde4
// cX,1(J=ANI>:45+Pe+TB-:9cPdd5CK;2S8]0\<g-c<c6(.?,+]cAOCY+5ZE,Q7RZ
// U34X@&WU^T2#JY)VJ=6ZMe\LC^H?IOTW#7PYWL2@]5C/0<-36/R/)T2I\>M@/L;-
// NA7:WC@d>g^^8FYLGeL]QJ9S6<JUNQZ#N<5J^-ZT;6FJ&>^-##)\fM;gT+BF+KGR
// +U3.#=V29P?-A,C#W/FTQGVE<;NV^#LaU,XF5TaT+F:5F:dIgR_BB-dA-;]K)bP;
// 0505^U==1P7=)85e/F<5>FPNdgb+1R2J<T^0HKcQ.8T2HVWMJW)6HZT:PTX6;;#b
// d^1P(_6fJQQI<)WA<96MF_&7THaOc484BgNA4E=4ZMg=[.@,A4b/f6^R20=@NNcC
// ;0-5bF)Md2FJ,.N3&ZF/1V]A8g&2D?5N)aJV;1-7a5?c?JV#ALXT]DP[P,4cI::C
// c3]6KC[aJYc<H66E8;&[7O:6@=]_T8DB)E\_7F1Sce2U[4UO:^KA9-+.;()RbJ<f
// +FMFN4<63IY/O3,\ZZ&1A\KQ4-EKZ\Lb2GU5=W,Db)b<Ne)&\-UM7VNT0d]e(GJY
// X5T:),_E/\(^a<:>E4V[d+[XNNd>4>>8dL7eCY:ed>X:K0I;A:c^WGgJ^,8A95.M
// R@6eS[c:I7cP(8cY[?-?62bNM-6&.M93#+L0R>gD-#H,;NA+g0M=g4#KIG^N]UNC
// F-bQ6-Ud++VE5#gPK4dW3)#E5dHM1DAM?3O?3BX2D=)^38;?,aW5+E@Ia6<=.0P(
// cVTRC81(Ad6.bEe5a6aC_2G7MVLK@Q9SH>T4+70X_NbV;XW@L9./]INbOK]SRLc3
// 3&IZ4;T<,=gDP0^G6B8MX.>?&R;QA2J81+O<8@(a9>[(N+.S2_AAeg4R^Cg6cR#D
// ?\Q^[KW2c6A=SJ:S+(D/a=LQ+]ZW=3b9+1,E+;.LcM91R]QR@8V]+JFXSBH[MU:W
// HDQ?L^HDEF#SDHP^I(1U52LCGY0-9EQVZIOH1F&MQ;5;NYU\=>(I;/NK^=W.<XbV
// ([Q+WSH)+cUR@\4.)@EH(T@eQgR//\-N;0XC,7,DT.KcR2TdcO<OYZ[7+-)La]:@
// DYd@-?NF+(]34bC:I,\7_U:Ba+6P#K(=CXR9\[3)\/Z#MM^d\K<W=)T;^6S]b5HM
// ^YSX<T_f/Ka8gUM+/27GJDTEV]UW@NSW;_d#I2>)/FWF:D+C2X00QHXDb_g,(:PI
// 3=J&]K0CG@E9@cN/0gT(1-9K95dO_CZL-Vd#95D/bf-]F7QPH7PND\2)d\M=TR:g
// K-bg&L5;MbD:VGBS5KdRCbW;e#&QKSS>D_WQ);&;T\HLFbg-C--5^aD#?#^E.:/I
// ;\g32XK][6Z=R#F7d5UX-8JB5,GeeO[655;JW^c718XFGaWeRY?SBH5dF):]U[K-
// 8:E-6<[e7c,fE#_6eaN2V99N0-HcFHCcR^OQcRRCW9LEEg4C)QB@>+Ye=(Y4c=P.
// d@F+./2MJ.H.ZD(]]PDN0-Y,YdT@Te#Mb@)-4VQI2ZbgN#c(QJHF,dQ)N@MO>0e,
// L&/WX3^T045YU-:eM,6^<R58&E;Z6dMP3<>H\@7#Sa<a8P+-D.CICLP@?\(K4)gC
// ##5?H#A,>5A\Z99BDc+VT?UMW<&VXMMLBFEQ\a,?O6S:+@cKbBbWbXNaa.@ec__B
// 1c-=Y?892J&YBHOBK#1-?b[I9IfD9JI05#8_Ha(LM]^.B+#92_LYPAH]Z<\P@QMf
// 25g4\)cUJY#N,c+CMMDNGRSg3JP(XGCCZ6.5V4V72M8QCMXfcBF7B6EcUN-KLRgJ
// cIN(T[A<bE+TA&PZ\2bX.D+?FceT7cHDLAVZN<?6Jd)/,9Y#,0QJ2-ag:#;>,C_(
// ID;O0DY#]O#dGA7KVKUK=>,:bSg[MNOJG_ZA)X33CVD=#J.[gD_>WP4#ZYZ=1F8X
// [Qa<1=41dD[2-RZNP,95VJ,ZCT7AK0SZ3&>-O5=7H.CR_g4A##YZX/eV4P7\\-SU
// e2eFf-_aJNV=VAg,#.L=><Q9J+2]X=X1?MfUC;1EHa2VVM:?4Z/JX[SH#24S(),F
// J=[e/:NfB2?0IB,eI]IQ6>_57_<2a2CY_8d58#=M\aMW1QPL.RX#Ze\HD_]#A:+9
// U-B.0KUgeaFMe>:V@d@#L#C+-(5>,E&27P&MQ5LI7N84&?DP@.:1/&S=.>-ERE&7
// ;f@XX;#OgdXT+Rg7GKVAdB-XcBRJ.c1&I-XFe)YIgL[IN+a..\;RE&E=53Qeee=:
// RL_JY)\f2,E,7Rc;AQb#gA9J93;=D1]^C7;d?5XBKW8XV5\]W5;.>eN33\:3)0BX
// HbPW<>&2\<M.<Y@UcZGBZ0&B#^3)d/bffN\Y64-4Y0&/XP6,V>S,cFWFFB=SW3K-
// 0OP_JL;f7#EQB(1[4<HL_4)2+<))H=O_7cTP@3SX9=.YB2fR(\[75L.Vb64D4.P+
// XW#,]CaPR:).Rd/M-7P=_c/f6DNP&&O=B;EV]]8gTANN8GUJ2dPY2DD9L>@@VUJ\
// &XC_c\f#JW@H:+WK18(4E(UYQYXWf?)^:QGU:S5TJ?/:)8G,KU:g:X3-#XJUN0:g
// (9Q8Q6d;2F)aJ?]_\F(59<38OB\ECgc@EEZ)WROKAS;MO;E#EAS)bSBXFY&H]4(f
// CL8I]2.\J7gC3b)S[4\_1K?Dce-ZA1.M\Eff(IV(-[P8[aQd-^[ZRFI.-O.J>#F+
// LD3VVK-SW/88^9RMMS(4X><[:,JF?6@f+?##L+5b9V>Y/F5<N4Q\&G9.J6]L&FKF
// #e\USFF@P7AM6X[Z)]^,c8N^,E>U->OU:bY0,]?I443O+HV7HfEVHEfUAQf;B6,8
// KN+5P?[<c:<BaQKa&;36BJd;J#L)&5NY\28G82V[a9[G5>O^LU#X)Y.V[OZd5Raa
// 9g9?UgN1_E;WK=b07TA?=W-_N5aVE&f@(=L+(E)@/9Eb+]0K\Mg@[?YL=Y)3_Z1d
// K:ESZ,7R\bNU03f8(YMI<PLT+P..+E?:afC&\3#]+(:VRQPC3A;:@3;g?[6IE?-W
// ;ZOM:ZeX(^8A43geO^A+<S9gCRLfg8NBZQ6[)f9[-09?O5Y8b3Fc)b;GO[)3CG8&
// DB,,F\9S2DE+K/(#W^HK\.BPA#LSbg.DDad0[2Y^Nd@J=C548RI-WFLb,E,;OdT;
// N-()0843KEAGI43Q;LXc+S3VMX2_#=N8/BP?20)62d]02_E.7+(R#gdF/JKSDA39
// a>SaQZ9cQ_[VB_(c@4LOFL@^5deDJ0<^(=:AX7?_HV=dT(:PX?I@^NeJ0K]NM>7M
// 0LeEa>[IN;FEI?H?6e:d1H1gU^NcA]TeNOfQa<T9MVH(:R<TJ_J<58#_P;.)0N-G
// 28:+\;f8cWR6T4.8cC7,IJ]/aAQM=dY@^Q/[,9T;GUd_,<RBfPPGGgWOAY4^J5B0
// KF+E-g]?e[;DDV>5N?34]14c6A(S?DA5fO]g=bFdJFc>(NG\]a2<AQG0.:V2^2\7
// ]ca8;MgN\^N(P[e;7Y,Ac8NKK37+T:J\;3I1UBWf2L=7&HL1d-7Pc,P,=-/DG/VD
// @DA?HX8P9,XR3/1@+B&&ec5:+GafgPNTK3S=D5e?DLET4AF>]eLO)P#0QIe8Ec_9
// Gb]=YMWU7CUZ,>5XE@b&F^C0ZROV(\&_ZW;ND>03B<]JYX?L[4]<V]T&Ig=;ZJKS
// HBUaAMe1MYX,1fY(a1Qag/b?a,TX\S&aW3KTUKe;78V+Aa2EII-OPZ=1X(;BLXDf
// #2&eTNBc>BeXT<Bf]<Ff26ZQ1e=+8C46Q;A<bXC0aN\.D0W-<O5A4#&>3R?.C=BV
// g+b+>gI0c-7(>T:+4L1GCNRX8(:,/b#X^XUfZQK?B53,-AC+b5a:1PW3U-1?0OP3
// Xf8,#ZEH3W0WOPdW4[=>g6<&.(82H<]Vf8H8R[2&cF(Z.a2:0(:gX>,DL:_f^YOL
// R&8:99)<Rd);.<AVQ=C1BA=C87OEgdbD?#N(8U4=M^2,(&AGV&_Eg[66DH^V>ZL+
// .W]IZ/L&;g;A.RV>3XUE,82:Ga@MD&[OHP[&HS;MAAf,ODP<IN@#+_RC@2Y0Z:HK
// d2UK@=]\2#F3)#F/WIS-O8;^MJHbY^C=7[R2FQL<Q:9\1:YP-8VRaPN7?O__<AY&
// ]g,b4GX3C>aTU4.7&(U<e()SFW)2g9+J3S;0Y_7Id,d[PDR+Fc?aN@g=79>)NINP
// _LQ//Oc(8L[+dYaLRQE>YG>Rc2Z_2WY3\#E.5eG(H4.7(Y(-H:K;UNN@G45E+N]D
// 9Y9Fe6MUHZ=3:6,6T1\\5-0SBE:7D<;J9@B4GLTXKBP,D^M4NQ2HY=.g_VMA/J\a
// <)3d7HfgFO_MFM^g00?#UE_&4F=Q^Nd/^VLKI^H-.L#:HUJU7,2G(6>XE(@6gK7_
// :NIQ),7EP:)cUcC[&Ra[R3V;5,cNQf]X35B<\-P2H5/8;Q5-C67KJTM3S=aG&1OQ
// 9a<3;:B;RTcUNaG\@fDY?D4DZf[_KG<BI2]);(_O=#;LaB-=BU9II5ELZ4Ce4ObU
// [G)RccMBPX(,)H47:5EZB@_-d,bNECbRWYFc\#-P^I[ZVfR0_>E1]P]H9I3Fc@,-
// ,QGdbN\VV7HH^Le;2-6:gCC-Xgd6SJ/-<^)GP#<)#<F7WB>-B<K-R5&F^FOP1Q[?
// 6>9L1(8_.b]Ma:O;GE^>T<RGG\SU3J?,N[/4TPS&B<-ZW]:=B;N[\.1agPDX3X(_
// ?aPT]N(U&_[P7<d&f4Z2(bEeM?\;g/QI5)N^F45C,&O-fe0SeAT<1Gf?L639T#<C
// 92b/EA.VK]4=F+>B0=/6+8/W,2RC494\)#0PWL)YQ3PSFb#M_I5]84b5CFE&FdLe
// B<gdDK0C#aJTDS;G#JJ@#dc=9=e1T0(UfF+8b1V/OGI(c(A//Qa+\D5Tf0-;V)@&
// G>I\-8&[b)fDT6aG68\a46\G^V[HX=eZXG4EA73-f+L?YR1SEBF#]g;dM<:P+GTT
// bU<2?H>d<SIP+/++99DZ,P&\@=EA-_IDQ,_N^,VML#Ie3f.4Y7QW8g3.J36H?PAd
// 35E+Yg&LS=1VYTb\8A73H)80eVHVUCVea-7dV8FcQ02f3X9<XC7_H+QH&2JD79Q3
// a3T5O&dD0aG#[/NRW2Ug<)Y[MI^bN/NQP[WDJF;[U2C^<;]QEN?@2M5<079;CQ[Q
// &T(H9[YH#529>aLB8X?\.IQPLK1S<gA4Sb=./U;82\1fY>X&9UT;<2X/O^>04D6H
// ].M:OVWYdMA#.NQRX3PP0d16LQWCK]WT9\E4+(1:T<)Kf+)b]O5NKYRTa&>[S_d@
// (c:DGa6Y@/\]U8D?FfZ[)OE1:5^_@]KfLe^UVg(QfEB#aIE2[:KeE3W8Ib^A,149
// (=>TN4>8eE=dPWb4TQ9.:d<=84f4RZ)K=#,=aDM339[G<aQb70II8ZP]7+&922AF
// W(=#.F[217QHAR,MMFVKYU^f?#WO.d4+<;a243[Z<9QH=/85d?P8e+?\1RH#+1a#
// eT6Z=KNeQL;/\GFEA;__CA,Q^0Vg63+Y_fUY</da2K:LcVSW)LU,G^UfQSCH0BHU
// F7bJN(3YPU,10Y6GV^NO\T#HVT3.>2a2W[12\(&_NRL2YITC)[a#:,W[AK>::5G;
// X6\B=C+^)T6,e4SCV&Q7EOcgYZ9QY&4K2YC+bY+OP;.K+W]QQ;FDdQG76O41/T^_
// 0Y&2PKQZPEX<QR_b:-]&9BF_PIY.TN+YJ3CW(6WBBWUHEG[P?9NF_F3g3SE9gD7E
// ^3(I9a8P<7@(AQY+)T.T\U5;SWM5;7VS@:TYPS\dBfW;>M/)Vd,?2b@2>DC99HN^
// Be)?J=f]FQ?F_YT\a:\PGJZSINCE,d-\GMBS?4ZUa-?XAYR)?fQ77\7+EFBAYT>_
// bF3NX4W,c81H^\.2^Kg)R4VINfg92YPUc09c36d?gV?KAV1W?HV(Y[/(G3c@;.Z^
// ,UMS2:^EQXUgP]-H3)KNB&f&V-RTg?\:.,2O-0G__Xe=d+0.A8MO0aUS.?g(c4X0
// Zdb/\QR=GWc8gW:Og]<c.;g)b9LMED>Y].bEX=NgbUQ\]YM;9J91C-Vg>>-BWa8R
// =JF(2UeLN6S31Q<GLUcJOdD1EK)@BOE@0.]++a9LeF\]Y:g-SMS^;_HA3X2_MGEC
// Q)N3b>L^F/b^B7]4PL^2.d9SSJ2DR:>,ZaXdC?6(FKRgIZg@D@VBPJ11Z)>egZDV
// <,:,^1<O]W5>6RDd;C6ME3K/KBH]5b89/&Q<A9&1C(f:e7<fW7<D<b^K=CDHQ9M_
// @/gI#Ff=_OV##8R0F?:DZ@C=CSA^^/_W?a0c@0Y[A?>(FgC.]6OG#C-bLEN8<K?S
// 25N;0cJVTfgKb<V#e46LO>bJ-TcG2MI^bgBG<XF5[7X/TN\E6Ne]>N]B333<Y3/A
// ZA73^MC\S/-9#,=#D#>V6VN7;1[YP9L82NJ&0\;URZB?@PR]1SNKfR&>8.X:NF0+
// NTT4KGJ:1Y_cY;&GZg<N7aaaf.?TeA=0-<^\d,4G[0FV;8,c1X>Ccg(7ET)T+MD@
// fg</:+AU27<DXUFF-R^15VU#&SET>aI)2-5K90KXC#)TE5Sg0_f?^K_cK]:CX>TL
// LZG>SMc7_gVQ(]X&TY9b]PN4S\X^4g=OU2)J.RLbIX-_=aFX5;&7Q)GQ9?fNF/[\
// U8_9^Q\2aYSFZBV;e5d:1;K6:6EGL\a6SNLD+9==GPYNA?ZVBeVd(WZaWf[f6),V
// D+XKTXQ(,HDb.8PVdJ/?.T24.9?a/]OFFdU)\REgN\I1F[8ZPTF^8)Z;W=Q_:GLZ
// ?@RPO4KSNLgSS6f71/<KBKP2R3GScN6+>]E=BY_#5eJ)LT\<7)3?I3TC7.P4>4,S
// NQTSGI,-??;00ESADe(OPOEg>#8XdF5f;&:(6&G&1))U_#>&:&N);Q)ITF\3Z-XE
// LF89O((9/8Ab3>RV1GM](gH/K#=dX<dOF]NV[d&T,&.AA2BPHME9M>\,,TRJ2O_E
// SO/.&XBJf:@[[RRU-_3ZL[^DOX@gJ7:PQ7650C015bTXODXC3Fa?5Rc6c=JOO1<^
// Q<cKMHf\N:>cg,Q5>HO@E#,Y0.D]B<((b/X@eQ+/9-_F^^=]XN)K]VZ-Tf\f:\0e
// ?\6E.<[e7ZeI[Z)IB/<IBE8dbJYaBQc2\b]1=?05^H=WVfTYH(>U[M];4_FK3=\L
// Y7ETO&Da0I2TQS7QI):3\E=SU:AM3JVCf-&C-5:cd9SD.3;NdEZ4V\WG1_cF_#IH
// VN4YS)X8@EZI0B5:)0NgBB.37BB39cB=QF_&Q.P<F8&LAL97D:E51-<<?c+)P:54
// 47S63I)K##1JN;=?:@)b;c6[<UM#3SG4dVCaQ-RENXTE53I/)E-I#7(1BgH54^LW
// 6dSa6V7;;adCO:3;1f:9?216<V0S><OT<@g3^Y73_GZQ5;cT(S=CZUGf.8;(73I4
// 1J1PB.T(DHGg2Z@HR_ARedXM7MJ)We?=VcO>PS#:7?AP(,XPL03c7_^\E.YL98CD
// ,<ARB&OSKQf>0g?;V@CeDQ_5eb<YU2.4E,bBK>>fK6-X-.]>5KF2XPd&NOD8R3)Y
// O6PN64adfVaL,c1;gg]Q47C+?,f15gNNbd(UG&ea)BWWFb])_+HPN2bPL6S]+C6^
// -WLNa,(Z(1G7IOECgEPULY+[Dc.&Q?T3;f^^)W;0S5+ZEC</H4(KJN:aM9.ZE@/E
// ^4c+=O#c-g+2gIb;)3eScVg]PJT2;BJS]XD.)@/5K;XD?C,[:W32XB]4Z]L>af^:
// <E,S:Y-((Z.>D?A(V(WaX>fg,C\AIDC[PUU2_#0ZL/a=8DQ02^WNL&7UfP5Q+8]E
// .+[<g(#(C/:C&))cG4AMV7@A[J2HO/55F2cUII5#B1cS9(II<.>[SAS[Y2Sa#QAL
// ]G7MLKM7.WO4_2?5PZ)A2HV#:0]DM-5KB..99.O&_P(5H-=1M8,^-F#7A.&+T.+D
// fR0\a(L?&C4#_P(]+N--,&YEcISZ&FB-Le1+P2cHV7;SJZU?9dJ90>P-)YH5Y5,,
// S5:DL_BfV:.6@bA36?@[8A0aQd3#?0?W=QS9(Sa1C0FU#N8M,2AF;4J_P]GD13,1
// (A/dWdaRR-.(MeV:IWd2P24:[UW(MCH]+J)UEN3+K[XDBcO3Nd+cgU?]^8LC#G<^
// \@(4-BdN2Af)5^+:G0?@23IMB.6Q,A;1N-GS\T0V8W#YC5B5[7OK]G:ddW^D0Q+0
// AYfX7/e,>@,e9<D8<<N)4NPC>_0XM+gV?NR5-b<WPIPBaG6R9:HD>+gaM:b0Y)\^
// ?-9GNLX;d-U963+PbH.d^G2XBD8IO/Rc1ZcKGIMfe20+^\=,FM1S/g#A^E3e+H-C
// 6D?N#TS3b0Da5=LK.[QVW7c2U9LJK^gO4fX#PAOOX_F/VX0)B77K@N0ZP8AJ^Ng9
// d>)7=HW+,+ReMUD+@R9b;b\.V=eP2Q8LDX[&(]?5VaBfQafdRS/_(bG_dUK92(^T
// fZLT>4>Pg]2CV1BWYcg4,cCa=#6<K>Z^:((11VD@QFS)\-G;.,C2CU_@760G6#,]
// 2>/V4I1e\,&(H?::Y;OR9OE78Q6:M1/0W.3FSP(-[/,BHC5T0^&2]+1e[C6&JZ)?
// 3KIUH#CY#5F<Va^-E5P7cUWF]J=+)Ff83&@<d]eXB#W^d;DQE@[DE[OTZ/<T0.^a
// ),aJDf]<5\OP=fYaG7,EQL&>\WI4FTA=RIT3CW7XP[Q2;(?RBb]JL3d1N>(Z/6]+
// Q,B.K80.5^4(MIA2cVR/2Y##P&-:=\T,g5H.#1._2B][T,)I24N<;_>FARb&B1aW
// GQ]R4S[M409(HAWU-^^&+1\2^/7-0TR<fGR3fKL#JW1S>DP<=:2VZNfDeRV_2/F)
// _gTA)VD;<Oa(0DE5?;bYBPMWBX0HMFHH0+OfdW2&11+b5K[[O6@+[4BV1aF+SJ/7
// c@:ESdL28eW?2V:a:b5&W,\G0N^ROJ#^\@HCFV1d1]))?aSEERO^RCZMX#.@U\f4
// UC3JR@=JXd#b-KI_XH@VQUL53gg2WegSVXZab@b+Na<]<B4?WUY5V(N@VYC>eZ3:
// ]()6^cW?;>0^^/NMf_<7EEE(;U51Jfb@CI7PY_Sf8;J_8-fKME(b,?IW(8XO--E1
// ,V@c/UZ[Q9:M>N9Wb<9[g&Hd8dV=54X&#X[RH8Ag[B7c<;.Y?O\\3Ig//X=L5MDf
// F2R.aP.#-;0T2ZEH;KS>HX)3S-A>:EH&Y&?/3Z8_^6VDRKZOSc)bTHVY<IX(S8WA
// 7BWDV8=A:0K9::C:E/BKZ9FfRDB,0(M?V18F6434AC-QHW;0,J?3W)?fS\)EJMIC
// ^?PZCG?+#aF24c7cNETV[0IGb-6JV]-c_>(-.=VF^c]D\7?5HaAXEQ7BW2K2WVXY
// ;X(c(AVWS67^0.,;U>3SMEc6)\YKL,T>^d@Q6TF:8]^aG4Q2-<DHW:-(;88LY^f_
// 2#g2?36A/ZeKZM[]H-.HX@9_XDWMd)TRSRA(YA@O80YEJH#6eX-;U70<5d>5&W7#
// O:\@XH)a,1^<T3IDT&>>2^\BZQUe#]?76J)@/4^d.7F:N6\OYHXAf8^DNb.g^VJH
// e=OVC([JSaQ>E9gRD:C#W?<:Db0_4_G3Ld]]dTA#?-OY;VDDE[.W7d8\&)5SG<#E
// PRY[G#<CEO@#GGA[BOX,SeTQcF5._OQ\b&5\)3bM,3_QK)WIYdb<I[ASCVXe[K:<
// Y0/fP&HCIT-_LJJ2>#SMK^T\:GaU5MB7-@Z7Ie2M2+e2MW,(WY?La0gS4J_6)TM)
// B#GX@E/0\\::Lf5<QH9@ZVW;PWbGe#T4Z\(IDaBL4HF;Be(8a^Y;e_A1GIH_:;5H
// K1PBbf5EIAU.PTf4<65b06ACS.[eJPBbW.g&/>(Z\BNb:Jc:(QF4bPeJ&@88Q3-a
// S\]3,+W:ZgQPS=&3QM>LbN<=(P813_,L2&H)>:B]YQ_A-NV4P)R)@.fOdA9bCeXL
// RCH,VLEPEPUWEfB2N,QE?PN;&O;N<7RE7T#V5/=Q=-3WfV2UKc@,\G-]T@O:2D9;
// T[BB#G??>f:Q@9LYGOU)gF8/K7L9XZ4[B2]\f)9fb-Q1MEd8]/ZDW^S#AOOIeL/V
// @UH4Y5>0;D+CcKFDN\AY_OfNLZ20P,P]eK)b9B3K@^Q5e(e-M\[-fTHYU1Jc&5E>
// W-R#->@/g-U<31^FC3-Y9YKI_dA94=FFTJ_=/WXC&YIYFS3[ScDfRT3#69>0O)+I
// S7H.bOf9[0<6)K_=F(19V@fISETPL@]\OLRJ/c2V\a3MTZB&4)V587b1_G:PMUHg
// &#;VfQYZKB_+TV/V=;dLPQBHgCLEM1_c\K=1[QeCgcL.Y<,]aN=2g#9&?2dE(&&7
// AH2V&/>B=-VSAe)7;a35T9Dafa5;RdA=dV)SK8NXSIO;HN@5R_.(E\>7L11_:1(@
// =7L1VULKedA2RKcIK>O2c/\5]V&TNdOQ?1SIU(DJYaGNc-;TJ<0;B3IZI7eLH?4@
// d\TZcDb94Q^OW=eXML.Z<MB^?FR7C>FZ@0L,)6L;b]_2#CP>()<E4(DP0:b#If6(
// =[ILT4Y^C[9[YLa.>;E9#+D[A]K>QGgbX&W9[fZ=-)1UHT+^3\/C(I,MLf,U+,E#
// Ub(?d1f/C]HQSe29aEFA\&;CY&g(U.QG.T\fd8NU);aOf=#T,A;+9:_^TWGcQA00
// 5\TeW)?T[_Nd&+8YRKZQNdHPOK;XM)L>3=C[58Cg?,5FQ;E)Q/aPMfD<RJB2Kc/_
// #Wf/Ue^/A,7PedNDLX-.K]-#GE3,V&#S1QDE6J7L:TaT]cb4BQ;\XR(Z+NZ&SPC(
// KJVF:96bS8-XS7ZWS]\<LF_BL99Z0VDW&f/1a8J5Od^PALB3gC;?1K(SM(5I&O3C
// []0?4[PfB,+dMXUQG5<0/FbAHY46<_c?D9+:8>8b-6Gd-VUccZ5.b)b4(gECQ6^f
// HUPL;QfJ@@2#FZCQ7++=b+g:U3daHNW7XLb^=)bIDB:d3)DTR\f8>=fC[B^bJ?R]
// 0\IM4d[HE8034\D@aA#N;/b3@5W?9?5=;KZIeX^[8R2/55/W0:=EN/PN_+EB;Zf5
// ,e@V^.CfaVJP8E(UQEGfC.G\TPB/0U-JaL86D)?/SKF=dDN[f.dL5TVJFLL#c9Ce
// /8A3g:<]X5+Kf08>6#D3U,E6)</V_T)2L;M)Z+_]Z7E)fQRFeBagR,,&gR)A2[aL
// LMMU5],LR>C,1#@(\cDP4B&#M\a/\ZV0/BT@UH9PdM5c-0A(VY8]_OZW[dW\/XZa
// Ud-N/_)>I\1H<UZdFBJG.DX0Ka]D^&[SQZ59a<CM<M<Y[2ea6,P-0A81JLXTa#P0
// (Wb0\SP:(=7,:I:bE_1P&#+:0YCJP5,bC/B9^-<<-f0\gg32Q]6CeBWQ/G:Cda19
// baA&M=HJ408MN<>QeO\[IY45dT3B_6.FLK>eJ0?ISLag4-=M)?&L0V>aGYBg=JdI
// :LVZTX]e2^:(5,P9N0L8)J5<TIPM&g&8>^TKKJJMKSa6;4NG([?P1YPVM1\//R3L
// P_QK\[.-J]:M:Me33=?b9d^-\JUdGUKgJXbO&R<[dX)ZVbJ_??5T3SgOaG<7YTDL
// KSFf-P.4/-XU<X#6Z10DO_BN=g?+W,Tb=55FV@cM[RK?S^=SLC,Aa#-]].R,JN^7
// eO0YHK(3.2R]F3(Se,-S\B+D7HA1[7(1H,[O/6&5[=^G4IAZTC4P[P_,,]V4dY\<
// 3D;[bE:KVJ&:_HG7&(3818I-?K^+_;HS#G1.\cNDgHCe1ZWbNdf4I-<aWJNaL=7F
// W^.gYM9:+:K_^e_)Re27AYBXVJOC[3#^Wf2c5/[\Fe7GdH7J9&D)^(/KO(=]9&W-
// dYDOgf78P#S,+_UgB[S#2dAJ1e,_GI+^SI6_R3dK6e)(X7)J]T=38Ve/;5=WNJXa
// IZd:TXL53>a@]:Hf3LA7\P6&E:&c2ZT=GeG&b@#ee11UX.+3;f_?9<_[@Xa_HQ6B
// DePC:03[BMC;]&/2KN1FWbK:PMI)^aILO1e6G)QYVAVca:7I<6+Ae2dGGC(/8#PQ
// 5;V@HE).;DY9>=EU=B7GNZN^ULYg1\OJ##Y&^G240YV\_K]]NJL)gY+ENU=FZ#].
// ,BfgaBNe<KWS:,WTRH@;C[75eC=FZ^<36<SPTGdM0W2A?E/f.AB5gBK3[TU>;<Z]
// D569Sd#)5b.aFY4P8_-#DMD7>CWI[GD,V;2HK=e+(T8E[IM[>/42GMCPJRW5JfSf
// Ag&=>DIM4ecYL0,@4KKWKK8^-5J^D;[80^P7,XB:eTGE\f&CeZdO&BS6dYVRKZ]E
// QIb:O-@U.V^b4P<@CTg43+</19V=X]4Y\GQ)AKMP+L5F@68A;8UebDdB=C+C=#UK
// ]ZP8Fb?N0dS9d?TP9,Y;_ZP556-V0E9O+PIH4g?c?Ia3W633@B&7NYQgT^3&HT^,
// fS))/I-;fSQ85-1V<OD8RD?DLceK:[g[R,?\UX+BX\c<#U_&J>&D>8@eWfd;@J_J
// _W;[1b6M,F<=,dDgTf[FU0#6IY_8B@Y4B9S0.ZXQ,[6AecG]>Ef.3BY:[CPP,I<M
// :<bP_JOF-=TS6[9T@3V4e\fSb26d+YC(V:,B@#Q\\YIOH4-RUOL]dD70b_-=5&K3
// -=)CSb+/^6fIYGSE7b?Z:NIB99aJ;WJ:^1]1g3&O:AB]-GSBX>6GT3IG[OPN<RgT
// DW+0fG63\ee0.B<Z,+\2G6L&cF<[@bSg=DF1K68\86Q6LI=f0+89d354P7?e1a)#
// ;MPLLfE@4.+bBLX\DO03TA;[=N?;O8A3,S4T[::A11QQXP48@^D93SJN:O>cAENM
// 4fO8[TX.E<,A2Mb\]AbL+OPK9:W-&5I.:G;We;&,MSS2;#dS11dRg3J8.#T;@a>(
// PQ2#;6M#V0\]O?TP.S9+5)#6N-c99g6Y41G>dX9#0-9\1@IU?UZQTAFc^>,1RZ_U
// Jff,FM>[6f+.\_D=JfVWK#U9Cd)Q?H.B]U00@^1g32dW;MA)//[KP]6?(9X1LBSL
// D9FKa;)(H2RAWd-?,-+U=fJ0;Ug0CQ]/<_Q#c<NH7=E[;I<26>-K(8><aLS5HK5&
// I/08]V5>UF6?@4)dA=380eR&JGOI9Qa2?-H+5H_b@+]U8_;(RBB&?Q.&4C]10aR9
// V0QD6H>3BgcM_A10MAU6)6M2eGa/JOJSE&[K[G-K01A,g:K/)CWQ^WPC.D0a(.+)
// O:V7#+LbL^QFX=2XZOIO4]FfZU@G3@E_/UL<+/OdJ\>89[]Bc3P:3ee0X.C(1-=g
// [Yb],c/P.dD-MCGFKPFO9[EQ&S^c<W+gN#=eN>FIV.>_bG>&W>A_<-://>Z)1CO)
// ?N1N&,PdO/R6-U\?><<?2BB9LdaE@/SP1-8HP-I[:PVL[SdBK0dA<Z+Ocgc^.QSE
// aQO0c[]YKM&Y.57FD++d6R&(\Vd_9YL;S4^cL-<Q&[f9=JN5@>_]aJ6]T8ENgMH\
// .=>,2gXGK5TB[]VWNUg>g@W(ZLN\K0+a&39<Xe[BGXYBcf+5Wa+?:8f(I#OI^?+P
// @-9f9Ea5d91e:aF7OI<M(-M-2^R/S]d-^4<bdAE#e27>]U1;AZ=EUO2I#T9e/I5E
// 8P/0A7&B3/E4^a410c?3E-C]I1MWYO^;D@1;[VT7A7]&fgP;;:BP<^7^76[f&YK;
// 09KMW+VL?295^;Fd.66]:bW/^=2=9]6dAGXN_QX\SF-ET2=M^(4@6T66<5@f5d4[
// \9baY+S,g@ZX8@QcE8KOfNURY@Ge5KINR]]^(EdE^6XS)ZK2+R@dVREWN(6FNN(9
// gC;a6D:HI>TIAHJYda>#_<8&LFOVS4SI_PK3YG)V(T#RHf(XQ2,5?:4>c1T,9K);
// b3:L25(cd([?>L\^A_?6WTE,b+9e(Fd<EKM<MUX/??e&R1<^@Eg#2ODZ;RA&\gO9
// ]&]J-K43Cf:YJPHH222[Sa8[I-,PgL+H^7Je/E)3T4)[?.[X+S5336.X2aO/H)N_
// eB1N0J89(9Q#W^&_>7F3MJ(Q_O<FRg/-Bc-c;N4R72,:U;3SALS5gA)KV-NAa93K
// G&E^/37YDdCXL0](d(AR@1WTDAE=XHbG8^)--ff=O8#BJAf)<?M6YB6AO0@8?X?b
// LVVZH#V<2;;SSHP/\b(N-^7V>;=-KW9fWK/Qf/RaP#eP8R56F@KH23+(^U)58Eb;
// 2<<Z].4O)+?c_SR:+Z]6,X8SP:cE7Y8d3BP&<<SPg5Ua:.-6?UTLK_.68b4DgR+R
// _L?T1G<YJ(aZ<NJ?_c[YW8-?9=C9-IO,,8L;Td5OC@eJf;aO;78S#U1-J3?Q.2=S
// 9YLb;JUC>=][NZ<O&PXYQSaL+8I_.&WBcSfOU&OC4M=JUf[1+>RWICK:O:RDA_4g
// ;fB/Y^(IZAgD7DX^3=e0.0;)7HXCHX:eZe10P<IOOX>HDW?L^G>Ub:e#@T<+WK?6
// KP.V=B-((f@8Va9_4>^1PU1d5N<.ALS>XG7RZNSBVCNEIWB,R0N>NR\/^c<IK/.a
// HV7@L?/-=]50b?EWfTOX+LTdL/JOI)S4(\\^.#&?_0S#9SH@C6U.K[]S>&gRKUgZ
// gfVNd-4>e1/K_5@AMQEN;T2_^6\6Mf7X>D>]/(<DWaLI&YD^N3Ica&XBF^Q>TU5e
// T<@]<G2T-fAL<U.2?01JaE,GYSSND(9,>:JCTLa4.49P7Ld0)FT6OOUPCg@+)@)P
// a>W,PXE/3Z+=J]V+[KY@109\F,5;2GKPBWC]@(FYLB7@7Z@gR&/I4fgb=LWVUI]9
// W/IbadD_AOZ+fO,@aF3#,4OYS,;&QAZ(M66R-LKfM<(SUL\@4fVWY\;b;4,JdgD5
// 9O@>L=:a.R&ETN3]H#H._255W;U-JgJgO=fd//YRF9fAEObI#dc7MT5^88aPMJ>L
// ;?=0/4B9]\@P7NUH&^:?@R8H/W?O(CUIe_e-+)?##[H0BQ))908W&U)L<cFGS<IO
// <B];bcE.4-[@\++C_QNb5M/aCKcbK&7C>4&VX&ZF8R<0d,;beL/CHE:P-F=.DBIL
// =S7W/Be912A&?6;4BB:#H+,LBR78V+C3:<LTM6Vg+;RC^gJC6MC/KNJ@Q7=C)V5V
// I\?;E8;)_b]/4]fBU-N5Ic&#AIN\8Q,76PP9?5>6,(HZ_ZPF[J=Z^E6)9@Lfe9+G
// TDNML/JW:BRI,a?CQ\ZZ;<UN#M:<<>@bfC[BdW-M/4cRW.)>^8V9:<fSKZY^JOM0
// .VRK[d_9,U;QCITPG+b9CNV20))+6[RMcH1Z54#0]XPV6&,.6BVR_@&g8gU9R68g
// b3ICTR>fC)YL#]]Od\M(Re>6#gR.?CXBcJG2]&?W],MWP#NFDE?)];b;-6_Z9Qe1
// =\G<LTO,B2P/07GZ\VZ[.(CDJW/WVI:[K_9=gF6K8#9KR-W)+YWKed.M[Q<eTC@C
// IbEYdae(H?4:FZMVUZVSR/L\@a]W?8AV>AOf5??K]O/(f85,\>[L1aHUHD^bPfU4
// M:[a]9:K2X-O,TS-2,]:S;UB[C]-F\H21Xcd:&]0ge6CSG,6=8gRFH[aC[cb#4-J
// =f=-a_+dK[99<f]McWg#DK;Y?/;.a[GG3/.IUG/X+ZB,&I01_&;A-G^8FUXN6+Y@
// <fOXRA\bD;8K=&UMXR,e[7F[JDK>0S+/?ag\S8.bD5YVE_LFcVg?5-bKA]ZJ^cZU
// \PS/:T.A-4a==@4E<&+Ec0/5c;\MXdI2YSM1UT/D_O3;==);KT5=\4e;8SVHO1EQ
// &N373[e=7@3BEY>TFd@Ag,DJT-<8KB494)2Sgg,M8MJRJ&N-@O\bEb9CJR56?>)H
// @Nf7)N@(.5@eN>\f_@0^Kg)E-C2TZE:,BK,^ZUHf1OT_ZQTaPJ/ZE\&<+K<X+RT7
// =b5aK7#DW=OT[7fME_EJ7FK7R+4b&BU;]=)R^6JdE=1JN<Vc9ZM4da=LEFg#6CcZ
// aQ@dLVVgXV<=IJI8W9AU3E+8K0H6GM_E0-e9)9U;6Z1S&-K4VTS=[7Ta,ZEIQ?.g
// 5R?MW;>,PDM3P2(2@g&.EI?L8f5ZP.X(6d(]:IMC^\U9FLNR_@BF-U;<GM+4LXHF
// D#L1[4)HY).B<XEYW/CCYZZ8F6S8SA>L&/He.L>?A7SHd4OF5&+686[c(aGXfX.P
// FfLC=L0V^7RS)_41ETbWK(^7:S)62gJ@/=Z>8g/7;O@CdSY_Ab19,64EA^1[fS4X
// _SH-ZM_5^_cH>[@+,0>H@&4F2G^eccED#A^PbP>PTHV(MM:8?(\6;>ZMWJ=B\/.6
// CSF_L4&G@)df:5H<-f9PBY8+;K@Fa3<_XgT#A,f,bGRJUH,8b@:c;O:,Y_Nf)<8O
// QTce)G:GJ=.M=M@PM\6_5PTF>J_NJY[-#[9C:b]S(A@PcT[7b;9IGNOD)-:>P8X@
// KRU5J_]0.>@[KL?TJVC3FMT;3CN-L]D=F,A)<.GB>3E1<,=#F>157=H[UHgBSPY2
// >@D^efW92WBJE>WW?12\S.<,289d<@[=[fN]#/K_eDf@T3T1M#9\T#U,#B@[[F-<
// bEENRQ>F#.CG9=7H\^Of?;1+;1g8bQ;d.#67@QKYOE<&_97b@3LICOLXRUH=eY0K
// Wb8f:TNJ>eGZP[L0D+K9JX3TXR]].PU(MTIC.c>+U?_>ZU/FfFU^G@_V:aZLg&7X
// GO;AXHNd7?8Hc;_fH6D^UO>Mgb&fVM.]H,ZF)42+HY<fW[+H9Q.Qc6XG6=.XC...
// f)-QT3]E?aeB3BcaDAK+Va@GAYRbJU-NI01f?YW_G+W+a@43NI7@S6G0a3g7>PVT
// L?3>Y^bNTB[-HIbO4&Z+VE6:\cf195dOH+MRJ-+F+aVPJ/@=S,M[FFDFbUdH-Ua/
// -/MXUAQg)\S;1UG4XgJ>gd\dH[E]g9)eb-R)#c^YF_FA22GE:LGI#)NKbZA?L2@/
// VE[\[N(MCBf9NW9F7\5E,bX+C6V)?9W14SVJ@IQ5[FCVHHGW(^XPZ,6;<@;<(CXT
// ?,e_X,?/^4MDPHB_UJA7d][2MR7CbAM\Uf[TgXD+#aAAd=MLQPef^O061,GZ8(P_
// EYR>,1AFPde@/CVGPDc-7>#(9I+W@gW]=32XWB[:RMa9;)Z2]_N.KSR,]3#7/9^B
// gUT&U4XZOG>\:FdQJA7Wg=0)C42O[D0EP8+21d,\E5cd6U-<L5Z:a/N<5R+T):]\
// ZdRA:AeSHZF5]5FIAOR4.QNfIQ5,BJbE8S-W(E>E)=eA\D8c.[P?ADc,A1OS^)d&
// 977USNfC#B8+NADZX[Y=:@g?=9..AMX0X_E&#6[aNE[XdB\eMbL=gc\29+gK]Z0K
// [OIZPH--<F;6Z+#C0]XTg[07SOW=ALEM6IDF)e^bIXU8RSa=PcB@.E96EJTP8]LO
// U7[F2MM,;[e[.SNNZ?L+CB7](FWS:JWWFYgH^d[NXaI@Z,F:Fe?-,Z7#VAe,1K_T
// (K&\]+>^UUdSTaK5RTT_DBCY9(80@-F7I1R-U/^<L3/.0-TGbQX3Vf<9<Z<S?MCa
// b,W,5[&cec+DBbdI6Q<Cf0SW2e&O/gJa8K?,IM)C1c&ba2d9(SM/);#3[.+I6?5^
// gFSIXVOP9L13S<K;Mb?E]6+(BGJ.))9G.8FD:?a5__1dVEeTV&<2XZ[,JJ=1)=3(
// Z@G>Q#@YAKR=0#XMCb)TF(1@(PW4DB__BgH&GQe,^506CIB9_b[_Z^A_4.L24#1O
// )>88<=,+0(IV.K&V,O5#O?g7H=/?L-;1V_g:N5^:R:KH>=0;Jf_6CeRB?N>_+,DF
// 18>:UD>)O:aSS:HaLN4-eG/)-b3Z5&K.Ecf?-cG?KMa0-B17@_O8YB(gBdQfcRFJ
// E^<3N&O1c-S@6b#UWFV6C2N+43\ZG1g_=fJZEK?AY&8G>091D,gF)<?3MDFb^cBO
// 0P9>V.L+/P;I0Re>d.FXB.=KGLSeQ./_c0G4LXf)BL:N79)^99&&2VLUA/0KA8f1
// _)X6PJ]0O0DdG3.WFE2#N43BgdMC&CX\fG()Z6B-E5GaDR9=fTGYSVbCf>eZ#7UB
// ]_+0M.#cI:OR,8^NXW-8VQa6,SK1&WYV@G1VBQL30I3?6(0<F7_Mfe\CN,@dY_N;
// LU6@0#Q-];5^b19E3[;Rac?WN^^aGL@HVJ:BC;:?#>AF^U(eZ,D4>CLZ;/:?CT]A
// DaY\19#E73IC_R5S(Gf<PY8W03M_7#]4ZFG874=XIC^S^HG]T]Y@)@B6IY#)PB=R
// :5P,XPJ,[E9D[6BF]:5.]^_VY/XF8IP,05HCA@ggVG7VJE>G\+1R<CMPL+d<f,dG
// 0/U&-bLA6KL1c<cP]0/Af;eRFM@E.]Q29D+02Q<OJ.ILJAfbgEEa]d<_IfT=NPaL
// cJHb#ULI1ILDC=Jf;6KV5OI.26Ba0DGfMWLHd103K^e]0]eLg7<8M22M:aF?K<3_
// /74c]@(V9M674f^AE&Yd?<)J2G_3aA2F.[6D2bI67B99)75:LEeCK0>2g@_a0Z)[
// M6bJ;H9g/-]e(71Q>A_]ac/GXHgX]G0<,#>W15Tag0aD_(&^b)I##L9OH<dXRS\)
// \(:GLY#AAff<XKVXPJ;1G;X#)c#.<cP1a+5.RJKG(52b;Ufe#_G>fN[cJI_(BF4d
// 8CG+[@LCDecZ_XPGP5P(7<[5H\Z>M0<fZGEG>46B#BR/S,D4cU^ED1V+dJ2H/T&V
// W8Yb5M01>JZQPbe?D(Q6#d4R:ObIDQdLC&;MXLgd?_U8?FZc>cW^T+b9\Zcd?Y>[
// &_KC0g3RaDCRO8^A(>7B-8+?(g3F<_Tg0E)TK?:YP6/eVG=GJB?]GS2[AfN^D&W.
// 7?M?,R\P19HKERKe46:.;P<X9=;N(IK5EX1_V6Q]C/\7)8#]1gQP^gS<J105/9Z-
// GdSeQ+:=Wf@g]E;aQBG/S[:EZPXgKY?#+H0^3W9dR-JWR+cc7Ked?8Ie_c.@=>7J
// 1eg9&:/HX93:^bB>dcQIP3/KMPPN0L.Q([>MRgZJZ[#AI6L;GIW)cZGR?T-dgVZ1
// 9F+R)KcaJJR^@JLSNU/J>]QZ3V1L;fMg&TNMe1LIZX]dFWP?1=L^W=ENZAG&?d@&
// PP1#U,U0?bfLA1\N,25G3)F;a+#4f&Z@A6Z[(IK\GBIKF-3P3>;bD<;)AcBWUW@D
// 0&2U8XBNId@_S/0+>Q49O4&_(+\8P1RPbeMbS7L,?ZN=Z6FK69IS64b;NDMY7DBB
// +.)6RC(><P0GTec?P3>;&:2>&+Ob-BFOUBNed7f58N1c//c33eYG\eHQKb@L+d_W
// fg=4e\N4>97#I1QRXWB(>gZ2-]9&<AKJdc,fNP/\AW=3SLf#cW)O>f=)@(9cXHR.
// K73Lga7D>G/#/(TQQ-:]:C7AL:8f/Y@^8[>W2VZLBJ<SNbS+IgHf9:]-?D;4M_XN
// MK/g\6Y9A>&8??F_,G>1DgB-DQa7?.IFJX#?&c6O>52&g:4MAYO/(I1[G8a9R:_8
// 6LOX;)TB30?dLYK)Z4VGU/NUB\J.-3=XU+?#cS:a^A)RgCe:Ib>Z\7LQN8aRJ=YC
// 7;M(_gOZL9EYR?NLJbg>93Z4:R[?53>J[fD#Z:Ca+Q6NDK\.75LeY?#9Y20YX0T^
// 8L1PL8MaL@J9/)NI@+fD&_J&:ZSR2STLFEf:[=I)YZTb=GHd^HM8VXX^&&+)Kg3X
// V]dXNGG_^U-UHJODBOGdc/-Q/9F5WBA=:;^N.LDQN\@GYf;N+>FeS9&S9/;#-CFO
// eUg(87/?J<VbO7]a7_bYb.N]80OVK8Y^K&e:#9Y.P&=1a9@deZcb[O&F3-EOH5:=
// gUB1;4+Z,e/F/229(Q3=A9CL8IfHT38FY>PEfdRGYNLZd^JM]R>K>#SJ8fC\<&6?
// (<<WEER89eG[g3]).WSdOVbdfFMg,,3RJ\XSScY53BI-RQ0;3)2IQF#?.4Ob+E#b
// 8-S0gFdFP^#WSg_>4V<6BU>0dE_bC6^G>J4RL5?[/@<O&:9Y[5S]-,HD-XcVH>/H
// eUR7/#+,YS+gC9MFfa;5K.M=@DA&B;W>B+M#;DR3NDOGSOEUCc(VR45UFBT\:7[E
// de<e;g^B[M:[5)=O,N[e,.#]^AEWe)2JVCY3X519eR3M>&2U5A#TV+a6AS0VXJ@)
// ;cWHWX)RH<3gG,WcA/,?F2FDfKN/4YV?YLWLQ8(1FZeY)eUg)U_<N^a9FK^a[]c<
// 6FQN)OF:0;gg@V=ZU3bcbBd19OX,(5U]J[^>>f+aO<UZ;6:P<)IE_8&f[J&P]QBQ
// PHU0.(d<9W@K^E7_cdG?<3@gBQIQQ3LHaCQ=\Ve?&ZT)67.#[#e]H0TWYMRU#a2[
// MS#=N[>ag.U8.:C]:Gf3e.<(;<[a@gPf+Kb,STQ\Ib.c/LOS3;Kb9Q6XS;C;T>],
// JJ+D\,R@2Idf79]1WK>9GMXa/TTe[VZ=b6D=A];De:B]bQOC+)-9/4]DX:&dCSAT
// B3-;dNfb\_1DM=7DSWS^dM4.ba5JF<.S]&]]JaY2YYGDVee1ac+gBS9SKJC5ScA9
// =PUZD=1X6V^^0/9&IRTZKXB#B?MaQIJ>UO?B<.75E9=0J5502YMYR6.<b=_-69f>
// ZcSYCXVdARTXW(JHD5BWCD]HYSc+(fc\U+Y_+c-4f_SgD>0DS)Sf]SY4WD+I=P5Z
// ?A=#(=O2/d\E&M83=aSMA578B@T0>HBUJ-^-S,L^5#/bPXUP<2IG5^07F52XF87.
// R.6KY#3-KY7JW,E6E?+DNOGKA:1;eVa-#(ARg2+WWe?/_.GFRK],(T3UL4>5W+&S
// @?DC[&&^e2\S)IgeEF6;(WCCD,F)JE,Q__TUKP;OVG43S&#gHB_1)Q0-Mg-C]XGM
// LJ^I8;#5P20;9>8.:HM&_f9(8JZ^SEDT#U@b@E863DR(3/c5-eXEO6_f;S#8-PX(
// [)#ddcGW/>C/?]THZEJ5;BK00=(,WFE0LUeM(7_-fG=AI3F\He9GRT1/W6[4]Dd?
// ;TJ=(FceP.U(N20>_?1aF/CaW.5LO/1P>1Y0,KI8ZJL:/=34>;X=,USC)CGXag5L
// E0J:f3N(J:b\EbK/7d;L(-#;X2&TB.&Q6D0LOIVY:LP)(GdNSH6eLQe<T43ZfcGa
// S=)4g.WOE\JET-Z_-Lac,XD.9GHG?#L0+J\Veg<FW(=O:<U+;W25g\K5P#25a5+\
// =_Wa0;4gY1g0AJ6)=5-\(AM\,<9O)b0NO&ef/FV[0I(NT_Ba]FDRd#QJV+,M:Hg0
// >7YXS#O&d,1;]KRbe+_MXR=@-6PS:B3CX:@e(QM3O-CGTHWI^>7LQcRNO&QQ:]W)
// 9>^c(1]Cd?/YC]E2\V6OQW7BK55U(dQSgZ+>QCaBA4_M-]];6=0bfgf6dQ._^A&^
// -_GKCPGEE2E1H7&XM_-H3gWZTa7@Y59F[Z>EMZ<N&ZGPcM4/2ZPBYG:RSIJL:0Q(
// ]I<GH>@MQWNN,J-Ce,5OL+Y/TZ\O58W,dA?b(b;^dC)&Q:[/e>Kf3ZbLO@dc\390
// 78-eSf-[24.H2Ta_=Ne<,UX,d_TeDe-g]0AA(;@V;Dg[6X,N^CX4VD]<\AIb=P@M
// aN;\a_9\:TP-AKI_->TadeQV_EL\/XZ:,Z;15<Ce<g:G>YGLU-.a4IcNZ2C?dYI#
// BK33QF&gDB?PAYV8d0fWTa)K=B&MZ32+7IY^Y]Tg0;d3VPHSM/V#CDW&#M>0B;:L
// ZREP#13O/F\C&Nd(]X^HFIgVF_ES16I9_H^+aV;IDU0@87#bYLcC(b)&25_<S[JA
// A[S=Q,,-ZA&<-3S3];JO70UcW;GgGDE(3Q),.LMc1YaNEK?b4Ed_O,R\;B:9Y8U.
// T#X?f1-5L#f>RR+.8S[gNIQGfZM#g&^R8^NN])Oe:O0(f@U7C6A@Wg_658UHYIB\
// d\cEM]\:H_(J/RX4-?.1]Ub@69E(V]M[YOPD5ER11c2NY_OY\N[fda@+-GI<&UQ1
// 2.-/6[[>G#\K@[G5)L1^)3UaRcZKM&];W-:H>5^,f1:#B@4(CQ.;d^8K42AFZK;D
// M^PX:)^?,(&?PH;b,+gdC^U=XFPE?I2.J^bF=1e5C#-@(5AT/g&8K^eZ+Nf^Saea
// Ka#2Jd3P,4:-1H>NAVfg]&,c2K+H59IIE(Q#&X\gJ+c47#gLI4IM6DIVbG^<2,7)
// =DG3<&Gg^+/OY(5JE9XG3(=^a7SE-VIK&-&FEdBgU15UQ<e/a\J[_0&-VCO3+OOF
// JI31gW<>BO@:dPM[DLI5VPYJ+./gV?c\^[&;a7//P-<-+f,_:aA:I;gBAL\3R2(G
// /7E9ZEe=K[A_^U_I&a:Z.G4FWbEP+1Sd>GNTIGN,&2fTK\T<NGA7Q&efVUS8]d+Q
// W/B6CI&bfICaA,51K2^KRY,>/<bF_9XHM9]+G@..9(,>+>TFM::?KPI-D6MLY+b]
// )I06_&IEY_R>(/#034?e@^&GKLXGT\V,2e3:,S,6_W/Gd3YEgLb0^/#gUgV/=>:3
// H-Y\;92,X;3AcfLE-\]@TL#JS5\3:CD+Mf8/&RR##=;a1V)M&CWVg^YNYLMSGX-[
// 6f\<]:C)cc595>XP<6<N2HL3U&.)=7FOW3DP0.@>b<#b3[Z+g2=b(R,G7=a]E+B?
// >V2cJ]?<#BK_]B;Pc)g5GHV;gI9,9BM=6]EP=7&3H21K6;PJ8G2O067PD[5Y]5@.
// dGS/TY1f__@N>LS)EB0HPY+TF>E9IGFg]=aeOd<@9&YC7P>#6()D+KEWBg2+TZbP
// ZIa>Gg&aDb&>Yg(g.DX2JNWO]4</)DHI[Y.I\6<].E\E]@F&D3F-V]3W&#UN3K0&
// 8^4Z4C>TSROf_0WT-dYPdQIDWNCOH1&\bL==5C9He5RYM&CU]=UEV+a.b9=/\ZIK
// 8O9[.&(__6Yf)>^>JO^K/7M@LMIOM(E6CE,I@.4LED=Eb&fIfL)]44F6FeBI]e[Y
// GT)Uf]@FHY&\KXZ#HD^+0OIJ@2b_H_M#LMWH:MMHKPZQ8]fP,0,O6THYGUN]_NPD
// &cA2]:L?VNNV&Q1?/UR+M:_W.&M/X.Lb_V02KKe#CdO(TMEf2S2/0N7T,#F34HA:
// />D2dBVSS#fA?@d20(@IN@AXFc(CXXdD@JBdQe9JF?BURS)@?]II0aa;7BDbaD)L
// Y3YO3FB#-R&0Z34J3DJ-(N6LAAE=2#-T7N42GBDA2c;DfIM_;?-ZQ&B8.,c>NHKN
// 4Zg:P.&A3I_LR[.KAI>?D]DP;AG0PVD200LA9]QHLV2[ES_18/=9<&U7)TPB,PEF
// :Q;3K_;5M_T/L@E6&J;?KK_W(L#^G#e/01=dgYcgN>;/_,;<??XMQ^S<?@c&d))E
// a@(>#V59R\DB^QY_J>?VDU+E7cF;Y509-;H,^,:\:#=[HLL7g(OG52B<JGQ._=\=
// _RCH^8F&L;0MAFE3D_-T0Rd=?[9e49f8S\WXYYLR9KH4[YPVG=95,/P0<@/d]6[L
// f7R;2=gMdR9c<c9ZcFF58M._?dJ;[Y6.EfG;E;.T>YebQ.#6GR213XXNPBSOYa2)
// HWL9;&F,\5+:f\d<G&LgRA,Ga71R>1^&YWTQd5;.;6E:VO>#SCDfL,P8N3eAc;J3
// HY+e3;AQNNLKWKY&MMB2d)+bK.eX)MaY-f31P^R@9/@9.9bFKPO<FdVZ6K1PRWaJ
// 1=_4-1ENR?O\[1>.fLFPX9IaQ]80>04F9[JM]2D=Y_#E\?5g(S^fM6ROD9@XQ^e(
// -AeW=HbI/;gG_0N?QIU?NEMWH4V_Y?V</+E_)N)RHe?\d]L.5@&<VgS(09D4b[,Y
// gcA/M&f,dQ1)feWK\a2Yd.CA9(S;YI)/ZK)9=e.ZKC77R4A<&ZY.U[NCOaJETH.O
// 2DL=c5+LgUYQ)d@\CBGfg^U&42=_=4P/Yf_U</A.I-]LVHFA[?-:9]_/5[L^9e+;
// 2//R<XFKP?[cSX5>gaRQ<<,A(,KPT:)X:;28=_0J7A<SQgYR:+8ZJT),<2GSF6eT
// 5b,?X14DT57dIGXK)Q;XgZ.dIKQfd19>KgB&Y0ga>-dIfFQOdPR1)J+_8S;JIM\/
// P_@>FJMC+R<]J]@BO;3)eF]caOfV,:56&\)^3fTW8D[Y_MGDc(4da#c--/F\b,Ae
// L6(DcBHFd#eU^XUJb\BD4>(UIA3JP(a)K4L6?1fHH-#b1g(6ADS^RO98=&V6]7\^
// FTZfUL8e<+a7=LfPVV6(?SRO3/Jaa+c1KE,\5PREc+IR::+?:-XeSCSUFPJY;YV)
// (P;[[/?U3X:8:(^Q,[.4P9[W_]94c/XJT]0XMf:GH?Fc6TNL0YgZf&RcD\B:413)
// ZJYJKC_YD)>J?33BB:/bI4\c.N6fcDR97dGBfVR3BQPe]OLTcO20>ZZ6C9Q7PU=.
// RVKOG=fQD&61DWO)ZN4Yb\R97e0+)=>F/^QQ;UK8K^);DQFBEgcB#Ld6ZW4[:-XP
// ,/)U=fU4>CF9bS<WWd/QAIZ?7P4BYFWC/3H=(QL/7:2>-XTV)P?-?6#FZc&,N>?:
// CV@7B:/.V3/2Vb8R-Gd+<,#\ZgJ]GPLCB819aO7D4.L012R[M<RE=2?N]0X@C:eE
// ?NKLb;M+3@KWU/PfI=R)dgdN_c-0f1gO-L/0M5H)L93(dZ5))eP.I,NLY6Uba8N8
// e:cZC3MP]=(EZOYIK;<WNQ2WZ>_:<3<=L.?#2KSPgNd6(1LG&fRULDdI;b-[T?,E
// D-C=<MWHQfLX@d-VI<3T9F^UgDF=Z6&V:@DQ@9T#A)bD:+e)QDd#N46@;SRG]Ia5
// d<B@.K:9)PNZ/<)-]Y0AH65aN\B2O8?X/Y&U6)E<@2L<YS(JFA-.915^M2I_d&Z#
// 5):fZUL#OZ[-F==X1d>D?D4+/C3N/8[(^BE\QIYL]WI)=W-J-SE0g8G#LD+7/0D7
// ]TYHb:6CRD6(CQZGeDSW+cM2d]F\3bd?FB\gG[IdCLRK&>T[B&]2[]Ma(IVGUEVS
// ^A-8L2>g4H9E\42Z2>#\_RdR&3LUX48O&6>-]RQAA>MVag[6E-K7IAYWLIWC1H0+
// .8TL95;[\2FHf.W#@<[36IFFMK4Ca\@13P5JD]f<-YD=<)^XTEZE<g>C1,#W.<;X
// ?C1-E.1QF:>I1-H12R+C5S0)H;L_-\R9B+g#)3,E,@<RCKJL_5A+BXN<6O]J_OZU
// 0?#H:7&FgNQdXb3)3A0M7cg2?#PBOL89eHF-<KMKU+D.A&>J83Rb6A@U-aG;84cX
// R>,#@&:d]a=bMfN7XM](TXO1E4BEgX=cONHOEg5N8W^Aac9QJQ3U)[OYLHa^OSFA
// >3H.IA@0[ZbV1^:MgJP2\U@UK;TK[8FB64S)1X0bgT+N<NRK[f<dPgDc1=GI1]5V
// 1>b-McG+fJfHAET,Z2FL+bFD&EAdESLWT>]bT92LU^;B4&QZeWR(Z(:7VdV=edBK
// ENK]I&cRHObUMI7X57^DS@#0XNa[_F;H>C1IaKO>AGE\GG[;7^>FBbQ7KY7Z??TF
// TA(]\A(-D3O)<XIR\:(;LBEO(1A5=O5S8O2PU6f2&a3P-+f.XAOgaNaJ,Q17-G4_
// RaQKB&@3Kd#=)-BBK9Ee_^Yd+Q<-B><+b0LH#]/8d\R8].7Ed_e1PVB;YZaG,<V2
// +F=>^a\F>?g7G#(R?Ua&C8T.KUX_<-IV2DQK_<K0GS@S4@JaO;N+BRKW<3Ve_;01
// ^6McJ)a09AE7.,KDQ@&K2\^VZdIc9RYC#L4-eD7S(6ee/BWE8\&GZIYJM4CT1LRL
// f;<6Ve#>NeFX,@+YHeOQLZfB(&7-PPB075/80>N-fbA\;,S:F65JJQddD\B\e,[O
// (U3a10Y^[cUCLO60I0LRR#4^a+[:K;10E/7Z,L#OMBg4UG>^FG5eY13(::C.c32e
// [IV.)a^T@VL\Y-#@QJ.)8@APQ.G0L\_8:G>4AV<1/WZT:b<9HHGO=9:O_1;-R1>\
// 6@f&,E;\Ya_EVd3^OR3P;^a#G7M@WIW,(aNb?FT+TP8Z@[GM.</)PULe[:bbE_a9
// ^K252e>G_8L+QFLJ7BF,SP>FNQO,92g)J:U(H_T/>7=7bI.0-C=F2He)OU)/]=^5
// (/6WadH)bF6Z;]YE)@35?;W_[T)4WgW)C>^O]?VW9T?G5QAgV\.CZg;IK=6?4bC2
// >DE]]/DT.9Z7RI1#O[VF@&fS4]-c?A.3AM>X6ZXJ+9Ne)Z0Y-.]9S-ZG#e,#QC/1
// T,EZJ.aS@3=dC55<9]U_4ODYBW5=\+C?8Wb[/9[AVIbR<f8=f6@7e4CW#gXcLg94
// 6#>D#S#O)FHGbd(9E7=[7f3XSXV/2R]69J1cQNI0\CW-gO0S69eV/-8[Y[fe-3J&
// G3]a&^H57@TI@d3U/a5fLG_-^g#[FF6Sae<[.JCf/Q\-&_gbO6IgSTEaKb84ge=D
// JAcM#-([5eQ]0Q:U.6EE0H:06>ILG86EN/KY/Y+I^DB]72IG]fDI0E;2g3-;32VM
// +7J?8KFg+S5dLFOW,0LW8_C.79H]4U0FgP:EN[==^M)9aS3P5=;^<YT_=4>9BeOM
// (..E-IE#]5^L>1D;C0E;.@=\A(<YCJ]3X/49],=/V<f&BR0C2H[^&B.S6KT5HIg[
// \+3Z\&IaB[_0<e8=>=/2H;F)#3VESG/#SIYc=MdcM9.H6]Cf0KfX?/MNAU:S\<:]
// ;ZWFXdA95\Q?_(U-HWb?S&,3S)K9T^C@ME^C;7ZZd/G]4f^PU>/)TYM<+=@OX_L3
// (&V/AFWH,3?(&<&]T.-E\I<G#TcdWWV]RT#7#@J)C:SI:@H2;&1)KR0.<&>^(e=0
// 9X(Z/[6\XA\a[G(B?FJ:eOQKNTRTA3\af><2/Sb#=?5K]+B?486Z0cM+N=R]3OTF
// @LHcEZMC/b9D1]N-]]gO2=7+dR73g[V5^N:](d]K_.EAa[&J5d][\2(#Re5GR)2g
// 0TW_KRfDVVSdgYU8CNG0KWKd#dC,@;3KGXOQa1(UdLdKbF^eg>^3e4N#TXTVFI7A
// :.F_8)LRE[GVQ)113N8<[<dO)+IRMB]72c9>gg,(\133AX(Z5=]E\O\MfM=HEAI0
// &BS]<S_G_Cg#X=WC8NO<QScNX>3]IQZ[7\PgbD_Ge4W_Hc7AaWJOA\+>E#FQ&=WH
// QVSNLR/Q2)aM6B2VNW=E.;<FIQI=HM[,G8,AegC-f5(3HN9+:(f7K]If^.Sf=C3T
// 9\CH^gEYY0H(FX\EbaA@FEK5AE>BJJ6Z9CL_LM-.(:eW+_662X?AS?5&/I?2bXcF
// b5@8\-.-V>C@67fcL(+207GSPDQgQb-3J,6NaKA?O51OF-KOEH--(X+-.TK2]PId
// 4:\2A>f/Y01\QJ=fCB<GX9.ffg3IJ,Ne/VTAc,fL:UF\[^?_M-XBL&+B@=V[HDL[
// fd?Ld7,GCU\cAN_U+-HdPQ3_SKQ_)A.WE+I1\Z>&CgQ,^ZbFZFX^)^Qc&b?gFWg^
// C@TSZM0C]_>SAgT,3FX(7DT<F1MdOcI1^9J9H.9Mf8BC1X55ec1]H@4A<EfV==2_
// b&c9?7&HX,0X(>aT2c3AG5BGI#A;WeV/Va_-gXK-XH9+-gS3Z5(CG]YDd8P1OE]7
// I?DY14>Y6\E>,?(,64d.Ub49B439&4:TYGgJ0RbQ)^F>c^<(U_BE;,NRVXCI4AIb
// YfaBbW@R\8A=V<2P2E8eP2SIZ_[&>UP8.1CXBE5XMf1-Y)ZBKHeW[_efQ\P@e9GB
// UI:6Wb^;O-T\1f=>g=M;g9K&OIP/,e?c[M,N.Cg:e3&/YAD2,F:\F8a?RT/0&@(U
// Xf_BP(@0]-4e+aU:I;dQM7N2>6]Z<K9<TB7O;^?--YN45^Hf0U3EH9bg\9AK48&b
// DQ;L^>T@K]F)Yfa41V#?,g7K.WV59SI1\S4847G>M+UR0OV4-]+6GD;?HGP7BC@3
// W)M6Eb1TT[(>XbQO0ba7#Cd0\=FL=b2:&U9a(31A/XVb(#;dU0>;2RB@EF]3f+[J
// ]Ab@cd)MM&)0IM5+GTA09dLaKX::SM&d77Q^QOE[DGL-0B1MU4e-DKd/^,?2:PI@
// J98FKW/@K9=M<@1=+?0RU5C.TV.fOO=I)RK.]CgQ<^/6U49bW^20dEI:P\O&):5Q
// =W(eW(H:[Hb0]X/ZO8:/9Q9e6a-8#;U/O^g6GAVb-KPG<B(=#He?.1-)H<ZF1OZ[
// OA\U56g0a87F6=07S<FK[WD\D#ME?#QeP85VMEGV01(dB[55SJ1V(Z)B/OGTe.D-
// #GJ9>9YC\>JI35#L6>P5Gdg1If7?QEL4LL8a1V=1E=S-g>4\2+=4,2[A?O^;@>dW
// 3K=4d9aEMDgAOF-4=3BJ?.GEe?#ZL;Xcf(aL[I,X)T(23R?C</=I.)LZ.Vf75eP>
// .g/]>3E,a>=<JBV-K8GfM>H4YgJ&QV[:1c2PYNUX(KedEGIR\&g;B8JR,)=b,JT,
// ]fcBNEaTBLKe.:&Y4/XUJLN#d=R9e]YZZJe4>:-ONZgBE,0J&R0[?0[0A-b1E^_)
// N7?M9](/5e.,VXPLe=ZOFK&Md=7BFJWJW(=E;=KM6[6?&;Bg3XK2AT;3(ff^BIZ0
// _MQRT^#,F0e)C:g^(8V/4<;GH-Ua:[0EXd^aef9@575A5KO33]6FMZT5(AGU&M[=
// ?7LN3/+V#_I=5#BD>S-OdYL)\[#,2Mb3f82\G7J)+Q\8@8T/J^7S6,FE+8-@.,f1
// GPKc^QJF<3(=2&5ZS_()O13?H?76:I.U6?M,JO3HGg)D-D]1/9\KQDC-bTE1XW;/
// ,?<JVP(RR0&#9U?/]W?3BD4]d1YNL+N[LP\Z2?5WYV:)RHPUAd/[3KI7P-NE5#a,
// cELJ1U@ZAIF99@Q;<K@S3Rc3O@c,-#W>1)]c5=CgH^Q#Z28K:?JGG5TC,ZU03>SI
// X+ZFLBHRD8OM7JBQ,35@?FBY09?98PXf-2g9@9^Rd;aaE3;2Y>P5X.8T)BPGJbYO
// >=O2:^_MA;U^NBC&Ub7gF]0>TZc[MSa1^J)/:]^GCQ]ZPS<4&(/3da6S@U++XYW1
// 7N[_)T54RO<\L^#:Q&gbABF\89SKU#K:)>1B#XVWH\-I3(V:<gA+f>D88YAR8_Lc
// VSJ<e4S6]4IT8a_^2SF_/f#Z(P<,[P&:8^5>;NL100^_]?f-UO<:A5X/2JdQXcI]
// F)(_[DXJ3I)C]Odc\cGQ124/PN51\OS<_(]01)@-/N.3H-A>V,O#\SEPH6L_^(=X
// 9V>1Lc+E/D&U\2Mf9Ubd+Z)JFdeGUb)OY8\SM/W1&YRCeLI;CZ+/>4DG><Mb1Z5(
// A-8ES6XAM1LYg]f86&AD6H^=ZS#&QT)g1A<&8.]d?dDQ,&Caf1<Y,>=-ITB<[&/#
// D#1Z=E]-_WM[&7-ND(Q=,X;^_EJAe0DaK^]NUM?F.HQS;XH]&^LJS?dKY?E/DQBZ
// [[9cOK)+M+>LTFEW34+&CcL7(U=[^H,QL5O<(L:A;PUW7;(d4(ZJ4YUMADN?=C<Q
// :O9C4W:ZA=\TEa4G[[@R?5I5BB-,8Q>4\Ef_=CDeaa3B),aZKD7_dbSOLV(^dE:F
// (Q<0]C4U<;US_Ba0R3P,^Xf<5O95,4(TL-@Q:<2@1Bc16)T++I/BbI4Q#eK]<T0R
// &[ZWU/MURVefAAR1c)RP>gY?A)#3ZXZ5=AE41D-L.ZFVN4Ib[5cP)07cI5.HcTD1
// =g81_3SM8)1#VQJBY<0(;+gNP:=1;C1S@R08H5+J9YZ@M&(3?=9Y&U.N:]M>K.e2
// ;E^?V.(_C=E2X;7-f>)=,TWH^M2dVOQ..;@QNZW@Ib[de3\QMCCU3+DIDaY3_\6O
// c@^C/3N;H.P^f_b<4[CT_ASbM,VK>D242M^T<T0JROM[fa7PF#gVdCMK&e&DH[2P
// 4#G:Q>d6-DY<62TGBQ-K07O(@Id48]dSUIN?DV8&PZ=/aY0CDf(Ye^G:U^)ga:XR
// U&7dP[-3ZRYTMMIK,.&3VKEYA.RgG6PO@];C6USf]eBGMJg@bEIATCd05]MgWNKK
// 8(7#Qc-Y9-W0>/=A78]R+E[f^+2K+e[YZ?0S=bZIbA;a_V=ca8O6ZMS=.;/aCUB_
// QT;4_(_e1\F?JOT.&P&=K?6P3b).TECW=&/F031@@ETfOI:XP)GY)^cF&NXbD:->
// >QO,9X-:,Lfg0EG6c==QJI[()TJC+9/DCgD_TUM2S]&H0<5,W\_ACKI@62U7(OXZ
// ,]3MPK3-d\cQ4e0dY=4Q6(PbS[ePLI>3OB#OD5<]Le(FA=TLcFJ/)/0DU#0b]J+c
// bF5U?E3eb^D+\..PB;5]a]f+)/c&7gAK)8NM6<-GFUG2A]]R+b8MR?AI95N7a\U\
// &-df3(cOP)L-,Vg-21AH5>6&5f8K>KNCLD(@#?14NY3A;?B2IXRMF-B&/6/>)LZ@
// Q6R>/I^1&,26R7:6RHbb)f(_KC,,LH89,-/2b1E^/4N5C?^2/81dgW>)=MDH9C1[
// OAI1MJ-#]Z+7Y5.Z@H]A&UX64.aZ(RdO4I;EO?BC4V\@N+OK\)<d2&AW-/L6Z-<K
// &9c++C7+<@C=,4>T.TRL+M7XHE#8CP_38eZ5NSa_NX\P2+BR7?df2MX0#\@)JK(7
// 574T2P6)?.YRg11b5.gV[6IRXcV#dUAN..)/L8Rec>a/_9e/7I6QRedUU0G7#9U=
// -Z__dUc^V#\LYM>gM8Y_U##=aF2e>A4SL^@JO]aBZKPVO_[TPRU<.gM.=\fG];d>
// FP?E[PU@TV5-,D#V)CF)597&OG)ag=#FGeD5-AGb:C?UGROID52ZZ=H]Q->-=YE,
// <;F&LKZXE9E()LF&AVA#N8T8SI;QWRK&2Y>QI-,T2PbHFEXZ[aRK;M/Cd&Y(T(BU
// Z6XNI3^SLD[9Jc6aN,CB#e5bHg::X6WZ1,WA9_QL:8b2:X\?/S49L@6K@?dE?R^2
// 1EgSM=YaJOL=T;XB#Y8M<I1OJ]<0LcE57_5TEL^0d0Wa=.FHg2MZ^4KFD/DQAPT\
// ?S+U0\^J.fTU?A2:d+7-C+^.X#7TbPX5c_3TG=)P+6WaGNHU=[O2HLM;(BfOd)6[
// -#2R[d8Z)=da?^-E4EeZYd22N?RVHF#,ZOHQJF-54aO]HR9\,aN=D=N:dCD@;O).
// Re7e8\fDK2c@aR5-<_H8FF/)&N-ON_W6d#d(>,8N146\QMRb2Uc)MZE=B,HCXL:6
// d7;5Wg?cXTGDM;D4b\K94(4Yb8M:aZF>eBAK)E.CEg))L/NRcYA+RC)4Y^-1@USf
// <QcMVY=Y,Z3J2J==f=Q8N3a)L>I]O<a0CK#\KNI;->_eF]+aVD9Q@N?OY#KF.^8&
// TJ&J8_fR<-F=WJ_B/EWV19VH]O0R@VNf5]?QDUHWcJgRVHJ[g9)a?#IMgW.#F_J=
// RL,N(A\.+H:Y[/KaP;fP#=I@6&aG#U6]KM6.fcH\(Ya0Yg.R]W/cA=a\NYAK6,,U
// <PVgED\S:=Wb0DJU)b7BgD8NbXG\_cVC@<#7[MR5.&D?cf23?c+NRUQ<aK+.Mgcc
// ?JaG-.ZBaa(/aD@@+Z/3_8:V?\AXD=];@[2<EJd&MYCFfH@N5]e+5AeV1:KNAf3=
// -FN-+WgE_PQX\(PX;RILW\22CZZT<T_T.SfW(G]=EKSD9>WWUYfb;T=gG-;@@a((
// [ULVgM1cOHIL==JFG1C:c-dUCcGCd&6X@\7\-^=<-aNC^.I,ZP@M@9B<f>2bfa<S
// C\E:9KH)3+YRP9D2aT^7V\CNRg):If/WLHV3V0-4]Sg.#P7&b5RHYOYV@;YO^F)[
// cQ)A0)?CQ,GJVAI15ZHDO9W\7GP?/=<&aEVY&1[AAJWgE-N[57[=BY,@:\07Kg&@
// (2LZ@N_c9:J)&C#1]A)ORYH1R#3Q1NgaQB6@f53aJMUAP[eR(&d3.[d]6UI8>WWY
// E:P;#4YU#GA+,GQ?+B_a:)a1J?YC<NI,83BD[YSX_J6>0f#[;#OTYa:fE=KKT\=#
// OP?KcaR_XU+-1f;006WIDf27616cIcJ,0(9F)ddbLI0+^G(7c__\C.M,d6>-TG8)
// K-C>0<DC;U<ec(WTEVISW2b]?(8cH[I^T[5:&FIaFR<+YbB[(\LWfQ@KG^P9\g]9
// ggB)0g70d&aE/aDK>c0<&ECfZW817(\<6IPQ[A2C_7KO=VA8RMTTR+I8]JPURc#D
// 1E5V7]F4f-D:DA]M(,6X0K\W??M54Y/OIb6@LO&MgbG\]CcK#G5=.5He?6+F:8H.
// &;d)>W/[M1d7H-ZXVH23.=EJJg1QDXI;83S)&=,W8_5Xb=K&B9Y5SR^gagM6eREP
// ,DKa)5,9@G51_GMf=cN3FCX\@WPN(7,=:=QcL9;;[#B7DC(JWNb4;7</-e6T@O8d
// BB-4V,,R[?RUO/CDa[/J/]QQc.]Ja3]K8T;V\]GGEeU47@D==#Vfe,U-6E>_DLCE
// 9WfFSPIW<CR5D)JH_RYWd_5D;@=@AC@W,&6&)J.2SJUcM74JJJ&K]cZ:TFV6g]OZ
// ][3JYUf2PR?DM[LGK#S::K@,O3)eQ]EI;A56/DW)P5OHAUJLHKD)c@WR9K.2^Oce
// \XQ)FY-@>;cAfCBNH>\A7Te[Q7&3\HXBPfZ68cb7;<Z+TO]VeM=P#YVa+R5HN)?T
// R_VQ\7b[CFALQNZb0.XJ@ddXc?;].T>7]7.1,T2FU/LO1O+KUTT5^LIMJ8?ABO4)
// (M>\C<7f73X@TZRNP,UC?,,(O_,EX,-T,?e8.D,040d)(HK.&8_fcOT6?J)gZQ(<
// JfRDe+K[4J?L3YG+G_V;I5Z^BSK==Jd.][<.U;#NKJWFBDceBb>c[X,4)LELK8>D
// KX6cMQ]^F??c;B,/2P_F_EA+I4?+K/E?@=:,@V)EJ\ZXAHLZ\KHN^?H#-ZIT==Y+
// EZ\U6,\U]1W9[NQICfaRcI:?];I,9b\R]=]&11,O#(2]::02Q+FP^Ce\>EGK1Y[a
// R#P([J:8;)BcC4F-R\ab6^7W-JI3Z9:A815/fN8D>+=4X:g-R<(+4_34&/@P6<S5
// McB<EQ((5WJ9(KWOR17eEV;^c6;U,;8]9\LJc(PbU>E+TSX\:6Ke2DfLT@9_YWF8
// M<cedD1SI=R.8&1X)OD8Q<4JbVGc5G;N[9T7fOA?fTZ_YL/2>8G3#NI4<M8:gUE9
// /H=XKM=XTZ+c^Wf^=J+[XKZc1C]g>2SAI?/b(;FAS+G:ILDB7O0M(\PFTL1aST(U
// RPR^5\Se9C+:Y_X>J>Z)24S93M?FVF7DP<\b79P>1>/]PC0Z5R?MU]_=(aT_D9TQ
// 9(;LI:@U1ZL2FTD(g#e=YBENKI,;/8cgJC7F6]e\c95N6_S+/eeG-DJa]Y])<V+K
// [ALb(e:Ld[99#?1#.??b,8:1D5fY,8<Rb7&c0-Q?7^SeI;f^:4U@O&JBT?#TD+Q;
// AI]L.cd+NdE29fIObYa4c\+/0Xg@?)EB?0_[Dc<+7[1Q>9L7G,0DH]4<D&LYbC\W
// 60Kf6;S+<ZgZUaXL0B]2L@Y[IA(bc@QWOca3+2K62<(gY1X&U:aeBY#M#9dVUGcg
// C(&,E71APT6N<dVSd2<Q/9UPHd/Y=FUFII[Z3)&gMTOUT4+97G>cE=PE]T_ab+[e
// O^C+XKgP^@Ib]SI6#N[5ZRZg,,1D==43(K0J-^JaEZQRDb@D0ZF25LDDM/60EB>B
// ,c+[Rd[HQG^g.8UJbO.W[BLE5f;(^:Q8d.b5(f@QJ5/gLaL9+:IBa;XPOKPNQ(#b
// WgG)KH]UA9478P-(ZV?O(.];0GQ[aF\C40XE(E[@JH]7-YI6T5aTO6eT,NIK5&CU
// Va[g;5VK>&J1?Q&B3Je1B]]cQ&cZc[_=6[E+=bHV1IYNLUR^YVYTVIgaLMQdYMcM
// )^7-Le_/2CC)FT:R1[^XFT50=dC5d]SOBV5:I2+</>M3VATI\L:>_IHT_R-Yc&c7
// eJ,7(Hea4T6NIgY]R&e2MbRPO)S;\=Y#(0N#KC[d,EQIXT[gP/^RHCe3>V>U<8M#
// ZB@;Ug6VY.8/.PMZC((K<L[]))76&\]=ZYAOS9KY)TDLX_/<]<egZcdC12&,a8PP
// EP@73UVWUO3Gc1=@<eNC=dM^YC3+441(CHCSG_Pd:aU,V2]9MX_:LFZNY2IGMHR#
// 71I;1W920@BHHFN@83AYVHLDR1d_<^(.QZ=c_YD/R_&_Y&A:+V(].15LDbWc/3I#
// 2.9W+\g\>5D8_JDTS&P8afeTVS0KHRZ;-[(@]=,1T3)g<TaG,C6@dU@:J7QTKNU3
// #MQKJPA9:@(-^<Q+AC6MS3cg?KL&Zb:^d@])HW]S0cJeFG:cg#:ZHQM\(//1[MbI
// XS=@&E,aLC7UNGBbg]72#XQP<92?UE=5-S:IA,Y8?PW3f:X/^)e?c#=T5I?)KDg1
// Yg#g2;;+PXDEPI=)WPG(1VP<_83OE]M#WPa^ZET+f6[e+KA9\+3.:\d3^N7fZc:.
// eNHa6?.:_<>FgV4GW79g+N6ad]IPMFCZ8Jf^N_^8JGDB?#JPMR?6U1eK?Ug+\_36
// WL;;Y;HY@T>dg57\#)W#(cIOSRd3?)3S4?Z&,>E1_B&\-](Y<9_\B)0UaLM>UF7P
// Ue<,6>#?M&[2CBZ6a<Fd&@Vb+TPM<E1A^X@;9e:H//).3GC66F7dbOb56CU#RJ9T
// -a]86X+OCI2&U.10;e7]ZS7:/5BeIWKEL^HJ5\4[Q+>^2Ea>DP-MAT(V)fccHT=<
// f]d4I-F?D_a[)4d.8aFe&7ZQ#dQRD:d.S\?JXO<?JcN2T[O1A1D]=BA7d;19R+HS
// d?3>]FH&U.F47d8SNa8Q=SFKFZKADa85;_PW;>=8@CUAb24YF6c&K:+GKG=HIF>W
// Z29ZZIa,9\7LIYUW=4W/;WD=ZQ7Z9(afZVJMbI51O\Hed+NV)E.5\fO;K>@KG@bJ
// =[6e,^FFKORQEg.OfUATZS]QIZY24HeHa\BeE+1GFJ+T1>D@TDLa,RIU/D=&b8NG
// D+@K2NL-6M/;DgdC00Rcg[ATL@=@06<g(@XKdBF=aN_#a^0dNc=@E=B2MMW1Z@7Q
// \.SS;.g[QcD>f558,(P6gfd@_2Q?^8NB]WOD[e>aM-ZfP#gY0U2Y))c=LI;D4W[V
// ?Mf4_S8e5D6KNM)70^9#4#XQ4757bTgV,eC4_P\A>/4@?bX01e6+=31b9K\#_#OB
// Df1:Qga;CCXQS-X[a]./37bbY)bP7#6F#NLeE1>&62fG8?3<(S@)NY&7[)=7-\RV
// SgZf3>M&__2D2YG6KN^CTaG2=.[PHU@e3IMLMR7XEN&;g&BMdY.[,4abX#@ZFHWK
// E0WJ=cESc\=O\4OIN:R99-D,9H53T)@L-PC-YG^Q]8;VJKE=SS,+7>X2E;YE?<-\
// K)_I?_b8PELN&Y.af2d,T@=Z,6)>JbMXb4V9ZaN_PKfS03d9>JB>,acDO&L&.1L:
// /R#GV,/]X[+3:>^=c6Be5>08Y1(7Y,WaTRRe7gPAKHaRF.C[WZ0TQ,[BB?W=JfRK
// 6]XX=Qc#7AR9;Qd097Y0J>D,+)g&1&UF@4d;Ic)42:)CBXXAe(=]6)#9&<=NfE=g
// CMa\3>bE9d^LK+J@YF9^#J;;ITY2\YJB0T[-.^fgQcI\:O.+_)I_]:8SfM@:/]C3
// JM11:Pc/HcT<,[G&1.9QMO]D[MYAY(.()?;Z3T2.2>04Ic7geE/dM2,#UQU0TOZ+
// aKdA,-\)_Z@S5HM&cJbM/5J5[96;9XB4B@cX,0ZO&H/fVfZTYK)WGGAE.EIS_I14
// +:/145L:Ya_>3&E.VN\J@X1fZ()-U48@PODGZ4H/53.UFPL[DF88[G#L1^D6OSJ:
// QFT57;dL>^;5C<C#bRBD:ZX+\8HIS@^/S(cWU1R,B(0gE^4?:5Z=U<V46@)#/;c>
// 7,I2]1gO;25\dR:E+5_3N9T3>[f-^A4<Z2@g]g^eUR64FLa4YMd33@K1+YEY_)<b
// dP0W&-H=C?,3B?=VA3BLXN3G^4Ug7DS)WRO6]9\GP:4J1a7aUGA+?fRJ84G:(NH[
// 9.?==8:3=a(YVM:@1=^..bCAD68CdHYLEWS4<TEd\F)(9Oa0L+LX[1eKUa78F&&H
// eS#A<6N\1;c:SCH#KJQT@[&\2I)NbX,dEg/CCd+J6@ZULV_)ES^Yg;?XO@PaL?U#
// G<+BI_R9WLGQ&ce_9\=U<+J:O=XQfAI9T<fG:+]K(URSNcG=gPJA079328,OfU,f
// XWPc7+:^-aU93@?d2@A/PaS05D/bCVgS?PRagPe>D6E]-SX:UK1&ARLY2(K#/dd+
// dDSa+KOHF-TIH49()_)S^M8MX/(G)=7H70(4=GdGB=:&R]Y;MgXNPXD9-ZQ#YF;I
// (#&,A:]Qb4#ED-L8APVF]JY=D^L:YaTeOW5W2CVG9GZ(5D5W#Te;\N]T\>bKM^=X
// 8PRDcKB2-USWK=&NOE3.LM@6N\f#0:/.b^4AR.RE47LAI5.C7.D=G@Y:BI[1HG[F
// +EMJ\S9(9EMK(2EXOFMEK8&2>HX2B8\<-(\bRccB&3JVUfIZ/;CZTXa#^aZ)#BTR
// 5J,1SW6VPKI4>QR3-Z[L>KWf11J.f9E.BVO+@GaIfGf>88/4RS?]7Y]8Q\Lf/GaB
// \b&O4R5f8DI><_AYTe>/(K(SI19U(3?c?9FS#eD/N,)3gTO,2P1ASYP=43<M)D#\
// U8I2#Dd>2a[^J2a+8^D@0YIKAQHXcOd=bJDf?a08CA<Z_25I5?@Pe^W4IbDAZWGZ
// SX8C4I]A]@2;GTRbD6\3X2RGYg2.&T^?ZS0XaI[Vb+6UCEe3Za+JS0>(,PMg<XM;
// <?,E6I88cLN3.+Q493[g7&1XG]VL8M.A=TFgdSBYIXGc4Og-L-]Db)2c/?17.Ga7
// bN2J/MI^7WC5_S47;:@fT)L<Qc28IfZH_JR8ZMd/@PJ2fJgaQ3cGHO0D]J_9C,VA
// I1WC#PZdASO/-=K;JL&:\NYDb;D?-6B1QeIaXM;U\?O.\bDg(bC03>cMXO47T3P9
// B(;WG\\e/[V,[+/)<#NAS#Ef)0G?2DPJZ@VL_f_4W,@UWFC\_X^?JW45\Ee02a-)
// R4\2QJ:=Me+^C</6K#&C[.[3<KXNJ4SJBBC&N&Y0C9gHHMe)Yd=-SJ[XHPYXeFN:
// EdNbMd<c_T-Q5-2+?[<DaA8=9G5Lb7;&644_(@<E#,3S+W-740)V_b?4,3R5XKbZ
// 9+M_Y1+0ZZTGJ+KU.gKcb325R/[G>1A(X>??#_D,+K<]9c9261.;],\ED[EQ)O]=
// eN=9f>A0(<MLAT\,F_4-f/GP9J2J?QC/:Aa?9Q_AOF\7>cNSGYC/ET/;O:,X6T=a
// 8+_MLL(;E0d9fd4L1_1.;Ad34Ec.UV+K3V4@VN0>T,M8WX/be1bH,[WB10a\41S9
// >;McEeSb+KHME,e7/5Xe5[)W,=\;TUG#AMHd<_\?3AHM1F0IdR.P&7U/JZb654<C
// ^,\0KF_;J#ZLf_.F6V:,e9d,86QYfHg.#HR&&gPU^VY^\?MTGQ@OTF/XIA[UG+?P
// 3EE,:Y?S\9bX\CD_TC7+bU\U3NTc7Kg06TfWDdX/VP8SV2JN2<HM5B?>5:3_R_(6
// >XODD1LGJ,9]D,B4WI=U5432Ug0J(e_@G@eH7QW?51b)QU3Y<,8\8_+3=fF:DJAF
// )U6&LY/)RQ+8Pe[P>/X_aD2^IC+fH(ECA^>HMZ#YK38F)f/(YaC?8DJB2D)0b/=?
// bPC7XBLNNERJ5GBP,7_e_DRL,E//CL<[0_26_Z#@ZQ?S;UaE<@TQ0H;&E_VWE-g&
// Ra3NO;e)YHJO8;BgVRe;DfWf?cNE6Y[K1-F?-?bV1KLIHH94X166+77P8&K78-YC
// d<QR:/=@T/GONIE-^DB/ATJJ]JB5(J9HO+[@LK#J7;GUKTI@.D.#+^RUPXUN/Xf&
// (:U?T)I7Y;dXSCFU4Q.AQcHZ2@<.a[HH4AFZFN/gQ2bP7WH3MD0ecf#5:>R>]/+g
// #G8+2OB9@9cM:Z?O6255c\FRdca717B;@V7+5^20:G86W8;NC.\g>Ld=(3WN@:^,
// QdV=O8>bVM(^W-]Q>(NEMK\5]S0[aPBPE/(YUDI&=8U^24GCXIS@SV?R<c\YAZ]O
// (Rb5UU&7f4CaT?0R.C67_c1_KbNJ&7W:VD?0,2@bUUJIY5D6EL)9e\-S#HEbCc;@
// [V8:9>;TZ+P(H1fFEPfH/N+YA=IFKf4@FL#[00e\PK4#AUQ)>?]ABY_82QH@@_TI
// &,=5EO@dP3eZ1)G:.OVWP,SEB35C\B;?E[4HBXb9DKLHR?P=)72[P2_(+g>59UU@
// Va7P0&85M2W;V]8Ie;AYEY#LY+\LaE#2EgMW&0Y;&OCHY8(?f_d_^/KF@[YPd>N9
// @VQ_6-ddeO:7<6A@]QL);4P5=^-)QcD.?)g+>6\LZPIM>T6.SB,7USXVAJ\(L?,G
// E109JBGHO:aTU96J](EI1>X40,cY@^UYA1ZFc_C:fX6cJ48a7H;U-90f65A2#UQG
// 4SR5S2/.F^>^OfOJ0(_^a[gYA7Z/:(M&?KH;DQOef9TN^f=QfK,PZ)B\:<N2:W:E
// dH64ZJ)T3D5[PQ2FQ4[;MCbg+#JO6(RdO(WK+P>(;/GR&UTMH;+HE<QPN1S7XR34
// <WRBcLNUE@4++09EdL7,<>1VEN4-93]cM4OP?8eK@)2f\:15-D0F<FOf,@BBM<fd
// )fP^.X5<TFPBPC&_WF(^8QS>O3B&f:Y6LI5Lag]&X,3dDPSZAcdOTdPFeWeCO<AJ
// 3EP?#eJNL_68?P5@\J;@1O_:7(COY>D8O+U4?R)0_E7dXc-&W64\O<#Se9=HUM.D
// 8;7YF0;1(Y;UPT?.?T.[4Ya3ILEQR<GR+,L@AMQ];>^_g?4T9cZ>/K0Od;GPS3TO
// F4ZgPR7IMY&<1O:X_SRI>:/(/6ffF8_[&G7bB2)GUg7TIeHQ(S/1W_=Y^?GfMYC7
// :b_-BO]aE?D=Z1C&<6+UMdM1FLd);]L;:IH367K@9PZ.H<ES2UIX+LR1M>E+E5g6
// HP5<Q.+O?)XN0N[Jf)F+8TeP=]U6)bF_T38a@;)XJ+4#AG1^?d#LDe2#3c+f+=Z@
// QO6,MJRT;9Y;KS-FQU;>G(=>45_PG?f2@N.GZ9-D1Q0e18&VE7.WX-+G\#M:]RJ;
// (2(UJ@DJ/+1Y8QcK#c&FK83UTP(9gP,d2^9GZ_?B@<YEg)e28UfQC0C5PD;9MFJ9
// <&X&F^?7VSAc#30XJe/-e:A7JcL4=+3ATU6Q3:\/[4#R<\M[F.Refa59eEg-OF?@
// +\O35-UNUa//J+-C6S_b\7G,7Yb@7.=b85Le0&AJ_QRWB8H0Jg.?4@IPRV&3A]\Y
// 13NQ;+.Nc?^1N^LS@g.)\S3bAc4D8J_0V+4C]W(:])fPQ#V@5\MSHUH\W8MEbfg;
// ]A5fe^TJ(:FD9gMgVM&-UM;KGd;&(GH)Qb#=_:T89F9K0<EH+?(4\d<e#4N]XGCI
// (_)c];<0caU<@K(]?JX;EPeU>=/T70XO\1g-1#E/a:Od,+L.>GPL4PIDJ+X,b7@(
// AHIE48?:)/N5T-P0MYI/7(e5^K?;Ud2ORB#W]/?O?<B##b9[Q_PRe)RRc9fPQWXS
// AC,Q/RV0V79(/&1e<0A3TOX1[e;a.VG)IJ8dBB21[3cF#EE-cQa,-4Gg;6D&,S5A
// R<1(5EXS;cf2>U-K005I6B55ZNg\;6;KJ-/A#RL,J53-b+Vg5f2I@:bR0EN_b#dJ
// A]FUL#ED@X/bBT-XRW4KYdg1C-NHF=(ND,,@8)7@5[I]=;^QDU.)>)W5,Q3Z;2]Q
// (HVG[?IX,cbE1OTE5?MP:7a90CWH+g2^E(4K7/Q7O=H)1X,&AMI6/3Y0:?OcSC5M
// U4Z=L6g(P#..UP9Ua#WJ7GII[MX1/F\-,8JL0ZCJ5cBD;5O^)O/ITUKWPZTG0H(K
// TVNS:R_4C1dKYZZ0[<cJ,Z<0QL7PF<g=AbL2=7e6[08Rg,X&XM:,]/cMcfc,8W4_
// 0^GZ.X..>OOJHP2+1\_5RUR_@-]<P]4CSH_@/aK7eX8K=992Z:G^.:;V>gHY^84Y
// 1V6;1P>][UUZ/,P7([Xf>=)@]6]>HP&?P/e-Aa/D)CU=/cSGNOb-IF\5#ZX:];H(
// T+YZJg&2Q#)gKdL1V;U50X@OQ4C^5#0R<c3@c:1d#[C2cdgI(U_MX2Se+J&5WNIM
// I>KB>K(96-95KEF2).S:068H_0?Ua/F>XG8GVdA)?SW[BV\=Xb7]MFO_?TD1gYBJ
// /b_D4,(?0W?0)Xc]_/H.>:X3[U]-_)XeCQ#I@&5B.=_?\5Z;JgaS<YC68W<KS>f)
// HSbLa<Za.>;:\MU;XATZMR=ZHc:V[OQFeFg&4BDZU8]FT4)=.(SSPf-e:\OUW0eA
// /7S+[5[+V;g.D)]]/>D<[bJEP_C6LfTPUZX2OKML57_/0Q-&:PM>7]+b5>8e8H&-
// \-K_aUfb=P=M#D[_gSb;JdJXGc@1#[T_V;+3aS9LWgP99IF<OPH<,PMIJPUV4MGW
// SE@\0\UgRE4/M0H^F)@N9V]KS#/KfP#aA>PW0M)_8d-T[d+.-(b<7AO\\[GJ,P/3
// \-C,S5g5MQRC1B4X-6F]HMX&@CX#g?K<F>2+GPA+QHc2<VF8EEIR[6140@Ibce2X
// d7-cCGYd;fJ4ED=[PNRaHJad,#6dgAV(fXgSG)@g,\^OM?&1VL1[T,CD>>Og&3:4
// A[5.+:G.6F-_L#UR2B8eX-MWUB5TVb86J9+I?UT[a+N0)-^6+56c0ZdQ^0#)Y0Z:
// gYe3AFW(&g<e\gD_UOf:=A]&C>e_-0[VZA)/##C2GQ^C4Mf\T\.#6U3A4b4f-UTZ
// L4Jc.BLZ2KN#_M)WBN25></].c5>4c-79Z(9a&&J;PB:J,3e;5]/E8978HK3W.6d
// 4(0,8WFVDga1c&&QCONZ@]Z.c,F;(Fc/T([_9-A?fe1PY@aMac9A&<ME-ISIUB9<
// C/cX6e\DWC)5@.(3g3L_(C69+eF83[]X8,I6LZ;d+N)HMQUGd;,eM6_aRFRY\+;>
// (;HRTHAXBKOU@bK3-UV>cXOVWQM/.0=;23]#[a3VX5LBKKX]@B9D)Cc?dVH9Ofe-
// fWW2KNeIQ](@?5D.S/_/;dNR<Ebfe3KY@P7(LXeE/4X;UD>d].Ag3P/D2?V>CS;5
// MNVO]DAO#2a:DJ&0+1B=EfC-+1BX4?Ab@gE)V/]]#N.WUQ,b(ZV:c\)?9J^C8_M(
// A/5R:OLT,@433.N>d]1@DVbX-O^0EJ/8?da[/TV<FKPSBb#NeZU^B82,_M5LNHH5
// d3&=&:c9?[A;O[F5W1N<?6Zb)2884be9+Y]GYc=[]g\f.TcM=g\1^-Lf^-I.(:e0
// VI7JDHPEPJ5Rf:+5FJYc3FaBf#8fGB9cQSJ9YW62C^<IBDJ@<>_Z7[8JC^YUN[.I
// WJ2K#\((C9<.F4VQCcQ@3W<?-aOaD_J;_X//37,X=PW62Oac_C,;-,V<D5gB7K4W
// X3V<]HJK0LJD&_2#B@&MKJOSa>Q51J@)XJVf.+JSJ=dQ_Q^f&+H;>f)^D0V;LD.,
// S[G;2?W-c]#<3A([2?[g9:7cf(+)Q+9UF@+)\2.6]^7^4aF)C=BF#^W733PXLS@4
// ;UH,KZ8RSUeaUPSdI+=68/9c&B6&@fV:-J9gN9SH=GM0&3f_baWVbaNF-1B_cd/c
// FR)W0X6F8f_4<-)IH@0_b6/64Z<RL2Y=48JYQcF+(@28GH]KM=1)ZYU.0(.P#EC>
// ,d3[A80TGVQKWMc1bBOe2VJ1]KI-&D@G;c=TR#2WD15+=UI<bYLTI?I]NI\9?BTX
// =8_6[._FQ8)4,BO1,<G_ENaLbJd=R];PbS8_Id#6DQf)f(WWcUb67W^+:UQdG]72
// N/.,Fd^;,@b_1A+84\K3_bZ\a,cMf.dB([T:^8QGOUU2&OAYVOA?ZeYX86S-b54_
// Bc?Q/e@D>THRd?8&Nb+GHXa5FJNG936]Oea3+YF3YAY>E@?EF\JB,fJC]LN2EDTV
// >0F86=>E\6-g?a@DG_^ce9YA8<;N]/@T?UL?[2D,@7>]XcAbJ>\S^K3@O-W?;712
// JDS)T+RWVJW_^+MI8K\TcZLdZW7<5UM-Q)E&HGdP/-Y39MGD)H/054.?N0@5(-0g
// L6PCU7:<]?@/cH(9?DRV_W.@H)4JU#4d<K1@N0D)NJIH=DKP=,P]XK/-BZ2b^@RG
// .R9KK<VTR=.IeJK)3b#A@[McLf]H]_3;VW8Ya,F98fG>=LMZO?eddd\?-bH84IN^
// Sc[PBG/Y.Fe^5T\+)bT(:F;K&_D+.,52-@NJ19<3;&a?EUKbX5Gg18GB.VO5A-c2
// URT]X(F##G#2H9J:5/B_Q5UCT^;X#aJHQA(I\@[=fJX)P=9g33-HU=V4,W5.7(0b
// L8RaU)/PJ+I,J:8QOfVSGQ,#I+K>1T)RL?+bb^a1)9&&6,I(RAX</fQ=H:OR<JJ@
// <JL7/8&bD6L:GN5C@LGc9a6O2JLF#YRK.[3,^+T4\0>=V>^>>:01#aT_QG3DD5EF
// f^Eff-;JSJ6[/Ud:^PZV[UeBL/SGG3C/6c;G3RSG7O=:4]VT\\?[RMQM:eZNC(R)
// bT62RRa>&XSC\<;+3?>K:0aMXcZDM72,-Zd2@=HOJ)X9\<X^OP2Nd[KZ3QUDBUI+
// 8_^ZGfF^-=+.F<8P;850bgHH:5e_?,[#OKEV02Ra+eLJ.gP_T]WTBMX3(Z5-.Oaa
// F7-\&K2aA[FSCdCJ)&I@O=5M7c:SP7?fP;HH0fJ4A\;[FS,U#I?F0BN7HT6XS&I,
// @+[XG<_/(+6V6NOLPd@4Ig,9RO59+E,>+8H?YJAKdUeBP:F7P+##X?eH:J#UUcME
// 3)?JUS2HOOC]VUfV@TQPJ\,@bgfOJb^RAE5W,ccJVBALa#M.[-6B<C^Q1dUS,b&f
// E&PH?P[,;Y?XRVdU\eDMWJJG6(?\.UFX(C>D(HDP>F=;@31/XZRTZ6C2<G6R</0F
// -BTG6KRU+A;7_B_6Y2cAXKF].7DXMCYa0]f\G7db@eKG8ULZLV2-c#NZ/c5eED\4
// Q2_(YK4B/3TLU?5G_.Ne=#_HA)5XFQ5CZ1,27-#JO+,W58bA3(<_8e)MTG.Q)&#e
// F3LN-e/c\a5[.BVP@K\H#U1FR-VD.][,M-Z7gMfM+,_JTR)De=UC_Y@KEfd(C^]E
// 8,_>TF?c7G(AD[0HG:cDZY]B9XCN](>X(Z/C?8,AA/^S[7RgH#,WfIBK3bb(?f=C
// &aKFX78&I^ASOAP=3,8?@F06S4;DIWb4QI6Te3;<g0Bd7CVK]S0b#T)50U:#\U?T
// ./Z+J5dX+V?.AU(_Ief89+WGU7)[H:bd(8A\V^\/&VgW+R;+A7ec=&_5+1I^I=Y/
// 7&9/8U)NG5&6H]IMfGG5\JM3WFY,)AGcS7<<P@:PWeKf+<YL_#f-4K1?E@1FTI5C
// >28g@W<g:/Y1W&K9ZGV3XE@I?G>RB(\0:\)0NZHbJC]-D?)Y8IB8A^CE6[Ie0TbN
// 0=9c#/8?7P:&&V^8H-e3@54P>K<81L0+-H7_^Y;BCOOBb0RI;6Z@a^<ES1ZM1&)B
// YcWc)E_F0+>1;XP=fP>ZJ6aAVA:N1J@:K&a1e#KYSGdS^cYD80T9(K&Z5&)X[Oe=
// 8N>5[TJ\TIe]]CW-K947?:56],GN]^+Fa7Ig3ccVDg#dN\0B5Peg.V0_b+E.N0BY
// 2[:cX0H1[b<Tga1gD\KWYXUCHD0:Y^F(7ag0+d-N5&V)AO2>9<#TRfBd>VN3-V@9
// Hg;LYaTY_b5=@V@#TZ<AeL^F=O4Mc).YMb@+_2)5E^GB8I6T1=;UL2NdH-0&.fV[
// XI1N+X9dOYNU9RL7.,FILa[H_@2&,>_U<adWaJ\)9<?f^2&1<?[7-\8.E<I\XK/f
// \S[\9.MU>:&/&8&GG(;<@03J>JQ]RFK/7,V=N?Ob4H#Y6+)O-70cEO4g4(U@BMR<
// ^[POLFGaZO/eOJ(K>+\M+M/+[\7B,[C?>c/@;-5C4WN@F:fILEYN90&dDI+<bS3g
// XM_ECJ:45BNKO=fK9^)YJAF1.I,76RggDDV&<W:BgM))4Zg&AI+]Qe\G0B6f-162
// K>]7RMRD]T76C7LP6YfU/+Q.I7)4L?,9,KMJYKIUc=B/SR\4F.\F=cb/4D1P-K7J
// 7F_,NLQA@+]T5AR@A?EACfA881aV8D1J3+RAaP]Q#WM#G>3\MA4=3QAY#(L5]?K:
// 85FJXN=f:-Ag^:^.\?(2^5EX8f]J:,.YHec=L3\<>:O\#()H/52&GZ3]9Vc,aTM)
// K_SBg<d_(^U/S>&_[E>^3SJ/F-(UeODJMQ1@-+RK(+MCfHWd_@-38-8/@[AfF?7)
// W>QbMa7JFa.J,Z6O&/;KBE0+A\PQ;A=A2-MBA\[][PZQOCMXI<OA7Y[MScL/cdL+
// 3AeTMg/T]DXF@8gQ#/.K#J=eXPAO)77C>VHeb203WA43<TT^Z]8eKK^[b[<DXCU#
// e.KZW:-I:(_OagY0?8\S9F1dRVg3#AT/(O^\J\-?_+_29=Fc3?5/1#YY6eN]XWBO
// Z7H112JP#cJ/07e]A8UALd8E_XRS8LB]+f(\LQ3W:KK@cD]4H\TYW#(I2W,4T3DD
// :AU(KUH0_DcLJ+F-5B?L3V;K5Qc9+VF;.SVL_:Q(eXV(C)=#)#7#MJP=DX._cH4]
// ^DAHTM6fC_MBgfVcHZC,^GXbRL50gY;,Qa_K<Q#,F^VKD/3VP)?(TOcK.V1C@eQP
// :0a&=UaE8[8;.BVCN.@ab/9XE+V.ZXJKca;/EQfCfDDa06LN[_J-ZG_8T8B=>f7S
// 0_^A?@B7cbOIOQB+5gUW\Y+^3#gG_^ZaIf\82F?aa.a6V;=-D/?WEd3D8K23HSHE
// gF/@9458/&?4Z9)Q5<[B52-g<.#DRE.:/e._4Q;JP86Y[1)TY>)]d@>,dDIH4gY4
// )D<J-GV&dabGEW,<)SV-1+)VTYXJb&1b7JQSfYHE4YF7T/7X1[TTX+M8.D^^d:2Z
// P5P^M01P@TPSIC#acHPg84BW72DXMGM/G02LXE<>],HZ#d:L3b4a7WLDb?#)7a^[
// [g8aJZ&9].\K1OK:Mg4E>5>G>]1G7=H6c:g<V;-PXGa/#V0e&8Mf@F66a#]cY64O
// E\G+41dd1S&]:P3YD97@,f;/-LM)=6H5IWK(Z9<7IaNG&1\?F;XK5L;&CLWgC]@6
// eeG^_7?18>ASS7fES<DO<92c<2#FbQ8+?Y6_)BA/[XSLc0NK[)QOS,H=LG=fF#_3
// />c\4MLT&S9./da+#9.[MW#R<cIGgEK.YRY;KXeR0?^)IY\+4F?)ED]eZIeA8>9Q
// ^gGN4<2U>O;R_[E1C^O[1d/Fb.BA9:\7QN7RQaEKb&g6M#_B58,69S:JN,(-_067
// AN4TH<]FP<E[-8C?>]]7QY=BHeT7>a344#R_=eO7^_,@3X=?Bd&Z(_VF-H[7;P:O
// ROMXDd:W&Z516ga>\^2,g)Va,ZY<&T8BLO?[#&_3]H<@-7.2_cY;)RMcJ>:&fX>Z
// N8H23P3>=2I=_=7],H37]KReWf?,,^]e&@D+0;N(_JV]a]IaY(ZLdQY/2[IddNS)
// ?RfAVAc@bED.=Y[?Y41UN<cY2NW^4VV.:..g[9#ff.f2/OCKG>Z8SQdHC-<ceIX_
// T[047>aXA9B?-\YIaXV?O^P&fe(Ae;;C.f.T3M#Q(cB4A):>\[cMK?[--6U1;e@F
// Ff;d.&((0SeV]M:ZE<H)b:5^#DJ@3\HbK;@FXD/S_F)fGCU^DAXf&(L]NJ@4f;:)
// 5LX9B6GfSSWJ?BS;gdgKQ7IS;]P(Vb^:F>\H<W6V/S83FZLA8.)aA]FeU.-T[R26
// X.aXO^MIA(RI@?F1/4&a;aK4^LR4&4Df6-fcFf>D)eC]P:[\]H=,ZNA6c.T\UX=^
// 75>@-]N_Q).HHD:,NbgXA_<VM+:9TSWRCHNda6P]GLWe&]_@g.>f12/H9D8SS^QY
// #B&_ddgeU&&dW=c^[HaR&-EWV.aggTJ/,/A8EHG8>RZ0ZX.ZIMNR@ZU.01)g_^(b
// AR13cEeFK<ZU3(_P0HYeU>CB2JW^2,cN40_ISK89:0\#A:3Kg&+G68FZ>@,Q.QN?
// ]C6PfCbd:;U3eR7),>#9X:V=Ba4P,=C@VJeE[G5b+33D.IQ)8@Y]=_//Vc?QTb70
// cDdW6.6\2R6=O-J\#C)Qe3Z=.S)<ABO6.E:ESZ[F75@+5GT#g;(_Z:A08L<MKURZ
// 38I:e@:WXD&]5,7\>ORI+9E5[;e4Jd=[T)\E^,9))c\NF4.9>M[5_X8,5Hf4+02_
// 90fCYP<J,9D(W:S15ACbP:e-8#&3[K;ASO0MbfB_]PC+<g8=<?[-ZfFaCf7BM;:a
// I;+AfDBRbXU<Gd=?gP@b@ZO1dAcN@:?T>KGAR3@,0U>b<TFG[4,GQGFQZJI\+-C3
// Y3g;D3&>S_<0+#eV(W1_?d&>0FVe<IUd_O>G[OTQH[F8W2P9.1QBVB=\(g59VHRE
// 0FQXLCDC9HEW\Y]A@.acQ:M=^U.GKXa,cJ.6\PeaNAf2f9F_ab)(bGM/NK7/+)Ig
// 0Z>G&#-Db.>3Rc9,<4MHV;WGC3c&egME6]I)A>ELKS(e9MU?M(QfdYa(I,E50;A@
// BS(6\0<eHS#SGZBgPeXOZDdd<YfQ/J^,0?WQ_9X7L[d99?<3e/D(O:.g5GAA:K2E
// JX@Z\ES.?WA,]-a)#MMSHA@3M@fg\B>^(1FE7?YLU60[/bPYJY?D^)U4Y:Q9a0)A
// 2gTBd);H>+2[&77eWQW?B)9EQMXf.KZb)<7c5EIAJ20L+I0]_VG])M);>B-<VTOb
// =Z.L4[]</(]6\?<_(8bL5(dIECabPTJD/J5,BW2ZO7;-5R9;EI&PG>FTJ)&9;C,\
// I-I8^-B4\\bJ_W4L)M4fYcYf4B[RGAc\ZA6/741.#_@7@@Fc7UOOBS#Q.CgeB&Eg
// PRH.3Z5LQ0g\JPYg-HEa_J>cWXdJ:3Uc/G-Z/a.-VG9Q>8>R4?U]7>84JUQL(,H&
// Gd)Y.S)&aS]KeI1IL:#0;M3,Ed=_\8_WDc)8(#[^AUJ-U[75XG80Q6X5eZX8<WRF
// =U3LYX2&SS@I-<B];TY:WVReKC=?Bc_Q<KC/ZU\?69]3g#^cLd^P9cOQ6-^T1,A;
// =c<ORVHNI,_OPLfJcH6V]QdI5-&W/;ZV)=U^ZA5N=[O2AP8K8)L[+dFN<7]:Ub;4
// _1C]0WBaRfFE+[AOSgaaJUFV4F\L[(1R8G3e)aJY<aC1DbX)>LPIHU5S]>)T0?Gb
// 9F&fK1D19P&.PH+Sa1CEE);L26;9J4T:QD7^)S-5S\Q-XWbB?B(VC2N\FSRZEK3R
// 9/4d&F[Zc1(\Pc)WD]5_(^8\OB9T91ZF1U^Qf5_f)CG#@K-:XN3[C6SE,FW=H.AU
// 0>O&#\+.4?K>:4USA6c]XMaSBfa?->^J9g_gV.Y4ALf11bSJOI/cU3[L.?[7KdX+
// HfdQf\>c#6]^[\b-/>SVeGe,I63CAOT01Y]TK1]FBDV?fW_FH(\N4egQ:M2(PPLL
// 9.[7&LXCH/fNFNd;67XO,7b&>..f:N09]9b[dN^JLcTA;<^Z(IWC7eHdD,7(#FI#
// 9/:&FNV^[2]7161.IAg8S75:GT?S(?b/AV><3_2[PRQEYDb;:=3GDSP+:E,5HMP,
// ,H_>G[5-bR7288HDA;EGf(XcLL^Fa;7\L<d8N&+++/Le^DQg/48d-PgO(36;-:-9
// NEOeWGdfgSJd.@#SH\)2d90_SYG&W.;JYJ3]N0a6C7.Y&3.S/VQ4H?J+B5G+U>T9
// JIYRQQ@KX;CRb4ASYdBIS0YV&IaKS(DNX3JQUKQ-B8=-1M1?4\1[_9IB/?bNN]GL
// ,4]QeRJ\A0M@C3UIASSG6E=#/K5NM+KUR=gP,LP2P6.>]Vd6PPJ9B1/1cd<]A]+M
// gg4_QA8+Zc:6e\Ce+1Lab-4gSFeQ+6_(06/VP^g3@Q6O5RG:);e,K^K;B:[f>8Y1
// Eaa24[D(MfJD\WXMR5[B2(L[Qf_@C>c-]W9<XabE4Ka@9)ZeHC7bPOLTb>W/7f\8
// \(7N#?HRI1YOIZbB1cGMJ/C>Hd;.3-HA1/1(R2aHB^\+_/:f-:7XP(LTI$
// `endprotected


 